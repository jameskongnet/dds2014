`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cgXvaBdnS5l2JIszSvIpfH0UzlgZSFrePF9eYStbAB3SL4d7KTVA9CUFxihjVCd2
F537alrnctai23vG1/aNCVAJY4dEzWeqYsHZSC6PlclEIQqyzwpLKBuaYeh+wpE2
5+JYs80l2MaLYZPhBycqDvGcThRjaviviPUbhHSTK7CUW6f0twBPh8Z1+0e5y6LF
7fOJD2vKVb76vBQErjQvDQn/xKpoXYYxosGztz2NDyFmeW34BWZhO3C1uIkjuLW5
II2NUup5IqxUgIztj5F2flQsxACn0p2qfpOu1chk27wOsb7gP2JbcwbYms7dl/u+
LxDTg7S5tHtSVxCa8ODyTlmFTpspqCMZG5wBzN16bCPGnesnn6RzGx6/CbCr8Kmh
Zq5AvxFLIedUoVwW+OjB08goSATdxKvkWsR4cFt75++rdg/2krvf+opt9bIwCQev
D7KIfFKwUxVN3ltQlUQoZlMX1vOZzAGdAKslywMC7Iih4HCbYAh0fXrWiuLXNIMY
skajaWT+Rxgh3ENbXGRr+h/Hh43BlnPbse9Fyylrt25G6yy7mWoWcAKRaDEu06wi
NhoX3+j09m7+Vu3zPTBj6nmtijc9VdhOR4YIOgX45cKki0EVENn+bH4H2wW0WGQC
j3xUf/w9tb2NKDf2BzovivP6QD1Us+dDP4R9qia3JWqvZm2tUASks8EeKIYzd2hM
WndQxWYbIef6C3jdsyx9uGo8OjPTs8qQY0ByS7+WOW68ZKgis/NSIqOYdKRFw6sw
iS7Q+NJ45KNdBBZISU5fp6NG5jA1j8R5tbMOCkGC+7ct1D+frDBGWuh/H9K5mWPV
j3GrnKPPfI5ipCZNdcjFlgkj3M139LpXIKZI1jwlcv3V6jTtmRuF9TtShK+ct3qC
giQhTMvR8PAkH/A6LeuL66j2fa9Tra4DreFmksWsF6VxX5nkkNOBfMTQsJtorPTE
jf7VSk0AwRnpam1rqnq8zNydRFtEd7nrrbWCFrikYHJAMD3fT7q3KbzSlFbIDihC
zip/1hLsYBSlTfGd64agYgm146jn6xCJgZ7T9aYB8c1WzljLRHxeU0KCQHgVCVZq
AF7pxZf2JtxVVJHiJ63z9YqVuR5mmK8dE73m37aKMERqy1zqqaIsAmevKutkwreS
ZdoQmtDJ7insVkBT1DHAR1gZRO4eTNHx19VDgetzjM59g9pZ8FSUM5954OZIw0bp
ZQ/oCIjw7Why21rERmFPomZcSFU5MkS4gsvqwkB7An4OUJb6B/oZ0ySH9Y9LE2us
FklRhhJfuX/dOuYmAGMzBXF0jc7R8by8tNsp9Tl2WLviQCpm34iZXX8TioTM58WG
eNcc7MGaks6B1AbJb4CFketerZKsqhC9xItJ+4mNokdkZ8NKYqjPqHOTZNPyJd3/
swK7yTQYlctYXCiYjwdAaA==
`protect END_PROTECTED
