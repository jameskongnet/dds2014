`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YWokdEFMxaUk5tuEOBmzRxq9peeW9HDlzUFBj2cmpPeZb+s9hdGEMVYQyn+mmbuQ
/X1OK6GM69Oo/u05d7MVbrPBORtcHWNQtGaYv55bfWYRRiz3SG7jE74j9hUxgw+/
ANJs60fnQM0D1yG0y9eRyezw1N/dGn2aGgXe3dacm7Ibafdw5mZgcCviNbaC36gK
AEoaG1gsE6kkpF8RedRnsUpUFAx1qmNopMYxFcxHSx2WPeFZU1cLJpNIdusPMeKo
Bh4MGCByD9o3i4Z3H5AMasFytrkair84UuSbGMCnLeCX19epF6BzFG8zP7vZl42Y
DT2ke0ZEP+Jy9qSDaspeATOzltR9/3CgZO5zsztBRyA17sJ7H0SBLvQf2aJxri/p
gBbUrGEuN0qBNY5QrZiCTZQ72NlV8hnLM78tTMVdp6+Vbxsl6eeroHmh0VEjt+dy
xPpc2iGsGc0Dh3NvHiLrOioboDPsjjXa+DStRrGcncevgc2gIdSpB0VmcjZTDXk0
hNDgyyIvnuMPjVnHvvD/0bXkm2v9Obayrt67U3PHWoA9/sgnCIe0gohDTDVyEfOb
4+aGk20d6tFqXjdu8XsNhzwh7Jm+aXfiTKnyefK0bmKDjYBCzNQvEKqbq8/A2xUx
tpCzfxyJI/G20SnpJDEYcSvcXZ4/jGmiXOUBRLpcCOWh1IEZPEOhc3PeKN64/qbH
tsUgMGbuY1Qtcz2gymc9xdC8AkVGPQrY8jkCP8WdqMpZr8UWkOqOJ3STwTXhTSt0
mRyChSr05cSOyTI52BtAluKS929KNnDkkCk0Luw7hMzF/90z6pIzn1QJVlxa4wdC
ciWYyCYFt2JDobn9UdVW9GVkW5GiI2edVIMS684Zj8l2Zmjea74NdSBwIKP3kdLI
nbZ9RM3z8AdgOQ643+Ih9N3ot/VxNlhU/8poxm3kft0bk/JJ1mh1t1gVunVB6R84
0StbSGqoB4BElUDkKU4+7JHfIDVaTAKCyK++4teI6ffHkZOM3la9/mjBT4wrO6uS
zXj/SZUVEN5YrHAqlvFd856UyFNAY/l7cXbVaBTUr50Wp2xmEbON00ED/ATVl6//
BMdvg8hvRnxYCBLDfdCewzQ7pvRggKdn/CKjDLofUZXxjXbqHrNmZNujWA98Xevk
XNYsOrQLBeL7Te4W+wclnVLFdAQEFYcCt85l4DevcJmy7+NsBnXRRfFy/b5n24ns
NXGgQqeK9tTDIgQ1ku8QF2l6hqK5azE2WBOF55+LeHTmkzFrR7FSeUtezUn8Bshl
SxZvDIBNnISZnnagiXBkpjDFZplCwFo1iNa20MCjcwNYmGk9g+GW4n8g2XIpEqkf
wWfkq6tUsm+s/NjiTnhWXfaib+8kowswtETrW91HWGcghS3c0q9g7uqMvHqKP4wQ
BUal6NgAjQSP9WlFk3w+C+ANN0u58JidU/7J3b1PdBAYIWBof0hhn3tZn2FwGFb6
a7jHuzUo8fBSAGCvAlaD1Oa8gQJmX3XwMdjfuRzGuW2oE1FRApGGaJFcLjoni5gb
JQq/+spC59QFQswJaAFD7Cg6yXty4VGt9AEE8NTcpg1KJCkyHJZow7jIFveCF142
YjjQNyYF95/ZIUcSACZJMt9Q/giUDwt2+6VBX0391FINp+PbnUp1jhH+LWmJ1lMs
mYEuaArUYHjg9JZQ/b9q+l8yYEfF62unqL8/72kyWk/YNRLvnhhbSC+OmA5ZNSC+
ilAhmEEDhJ8AhS/gT9HW6FyhG2RWfOCpQ1CP3Z31C14fatbZUXbE/lTYdEnXnCPv
OOmCX535STjEjBlV18rNOOYu5O++z21jQBPCYZ7E6jqsfCudT/CUIxStNvt6ohGK
99fiGWbrq+x8henLIzz/KyryVai8cwVMPGZybXXPNs3ZHUn4wSQCzRbT3Ti2w/KR
WqR2nJN/42/dXXUZbqcsN/Q1MbE2BwkblOWNwjG0Xgs/4bMRIRTypzcRNi9r84A1
a10cKJhsKW9iLdI6t3mbBA==
`protect END_PROTECTED
