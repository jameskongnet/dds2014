`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WZ0OG1oftcn0Rgl2+g3BB/bUC5/l4eT1hpTbQIfR3pxA8/4xaFZXSVrUd8KC9RHQ
qvrVZb36O72CDRu+11WFyQyab05vmx/IbEPuXZ7K8ZEthyGKBRaLQFg7qeeOUWvA
PSrxuoze1b06QObUBBqURVvUdbRkJUt/dbrKoWKZCKZyfc7I0jeOwhwkry/dgxfQ
tx963Hp5yCWJbfQn0g6cNXtGUyYdeE5xL7V9s4LLoHyBw1QTydrH+ftra56/mT3U
W3XStennYZcBxcvDoNd5f5J6I8duIFGqiCRAptIMUV2uOyTIQ31rgHHbkVPyDWEV
skX1K92A3BpfyY9j9gZuSzLl3f7XS4AQmcuHctqPYbdTv/LzOR6tBmE2WqhRnqcq
SGaHVCBTL2DgQSAC5pzDXRww9hyBAWBnIKOKM0bfqb4vkL15qJl/G5l9EGDUiHrg
kpr+9h20GcBgbNPV4Dx0bXEFimnEnth0Ryhbh8/vyJaSJsXEXfTgt0O4G8kjdSCN
AhkAsvrq5VZQXDFvvH8bJlpwKIy+aH/KPPfo8Kornv2fFgvqkHNTwJhN8g/wF5kv
HcYI4Z7ijwomTufvYeb42HVVIZpZN/jJU2yOQj0iKo+mPqAA8U3tu+GdAH8myKnE
pitR10JlG3DkkNibUZLIDhi/2K1oANqxpYODWFgOjCMNIz0JOKMg1gHM5nifTS/1
M3JSqdGVMhJdWaL4jcbc3WwyU1rdn8pxNvaVH+/HdIQG5SFG/EJKuxsgO7xeh4oq
177PCsVxsKTcy2BJ675CDUxeq+qyXpyZcoteTFikxuUcrYF84BGXBNgnV7kRbGom
yZrrJpPyplcxy+G0WHFWO+smI0CXvHKL7kraUpgLfmhXhJprloOC03FHlZc/q7pI
nwKf4USOlNNT79TtPFgVKJaIul2VGFf6+lAJSRt2hj/nD6noNRczCxSQdT1XFyPr
6laSBOmjKX8iKdwKRPLVZ3zzBUuFQt9AMMeK84aX7nMNHTk9KwfRmmIw0DmspGK2
7lXHUryiFqGogxFyNeAAJQ/WFEpdKSYAkkF1L+YlPGO1r2qU/KLSpn3CN7T469Bf
vHsjYrUlVrQEQKYtmapvXBSBOkpq3lUqz+3dIRDBzjqRE6dPcLARfqZXsJeeiqLb
bnE/dWQex2/w0gRQO9pXqyZmVgN928kv1gu3zcUwmzkj1nyctayYcYdmOtTkyLHq
D9Gd5UuJbR8aV0sK8XUUuFmgE0/cQ8qE/a+544cdrEtx+d4xecCXs6X5ccKkEfXu
Vq0AcH1kXQXgGUv/kYNDyLn/XJ6EdRIBspyPMQOnhjiYyih2SoccVZ5iBF8FGWxN
bfk41lab5PwjrtGcnPoAQkWIyiN9B93cP+0gwWnLYzTJgFtlmA2v4r+eDA4DyvFV
ZUq2apIaekAG+Rn/Ef84AA7tIgIqmBAHxx1+drBgYTsDIuRS68j1g76B4w92aoAM
VfkeZQfwFfs053gsFkveMzZllOxnrRAHYJ8t2oxdfDZ/bY/BE6lBw+lnvoM9Yl+S
HxJ0Cyl4H1QgTfgpc4Jwuz+yTMiCk7ydrYqYC0Que1HQ2yFrBollUcCL8hiwzthu
tQwHWTTtCrQhRnQV78NvQr9UWkPuGL64ZytO7JGHh7iAd7SW3xjcv/9yk4+yDB7a
5MABUUxDQNJJAbstorsoLpYzs4M/H72WVmxEcYdeGJ+0Jp1y2PDRSnqks+bYJ2Av
Sj3PGP8mchAQ2OiZc7ZXAyolRJaY3KEss7mUvEaT/HYNBwpvf7PRt1kHKscpc+ww
BYUATlBEethRaj7E83B7MLP+3pHD5w236vhfGPVwYfp8Mx2Hustd+lrGwVdp8g2I
BdCKd+SQlB8iqnfcQSb+a4z7yhNP1Y8spvmOYxiIkYGTOSxldQRi8DJsaf3BOnYF
bsWc01aBzhedLgdaICgmqnpKEW3MhlNHHcKStbhSsfmh+CnBOUyChsuKa1wLqS5W
0aEK1+ZHCGxII1zisou+C2jhh25covHUNMYz/4lt3W9J1qvzu28ZsRo8GWTRYUc6
2HFX65jA3zOiWx/AuSmr1SeMOxuZSBRLF/JUGc3MfCnt2iwsrAgeT48g5U5QXvXd
EmRKHOSwLGVPAh6Onm3/myXrv9YiC/tiI+CGlMB9e8Q+DIPdknentluyFWB0OJmK
OrIW89bdi4be9FkHv1L18xjld6gw6SC81/Gx78zSIgk=
`protect END_PROTECTED
