`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WG2YtDjXtmGv0He57lV5Vkn+TdTwpQyFUrX3tXFDfOsfihkLjfdqCcttnIIJj1bl
A+OAvBa+9QF76sijeBVg9Fjru0524DNq6ISFlsuNASEFr66jmI2L00Q5Ztq6DinW
UbvdklzbxQlg4Ywbt78z405U2yJ8bjTC3cJUkGog1wczpTqi1ttHaYxudom20X/E
s8qQVLHBiJ0XIxGWCrRz0bETAKpx/wgGGrtweCEzkoAQzHC/5qztL5fXFJTUBt5v
RQW4r2KCvyH0+Q0K2exCIJS87M3BVcOYabhM9dZ6dmv5/iFrEWzkHSxfJiaBdy0M
doOv2Qe3BH60rAshlDlOeNP2+ZKLK05qMQuHttObElySF7t8NmuPa9JaR0PKp7R3
SdKYjUw8mcSdrOEFYVvENLvzdYH/qqppwRV8jKqe0rcHVXiP3oDkYMrVff/AYP5t
mxLrSpVQBdFbP+xcWHf9KlNsrxy35vYFdDwIZ/fhx9lxJdVp4t9QLMfQLMeijk3m
Dt1CItGbTlAQwlpWN4p3X7HO69xXjW8KqNMwxOchoMeQWJdh2l2onLFLH1GXfFoz
TZ6h5jjYGP2gR6LN4yVDJAUhFdIo51CA329Xd+28tPFulAWi0vRB428hdnnHHAty
r3uQ9QADrzl4h5gp8aY1hyI2rS8/9RVlTAwCohaUDy9XmjwWz/C/ala7EkKHUl9g
oLR8KyaWq1S91vDpr8Q1WR9GIYB0dpRT1H67SDWZi7aiqOJB7doI4hYiuTjgTqlp
LWATFdN8mjysCdKQJSI3sbIhf7T6wlV/nsagtkPkVEqkB1fOseNIOq1MIxCeo/av
dCIZeKGj//HsYfZpJBn6JedJpf/mSKau4gs9yh+bOHDcANH1AlELJAjYUnikWHGe
MoBEYHcnqc1fhRBi1/MluhhgiQXFxWHsT1grOPDKGIeaJrdHlI71SFhiDWtR5sTT
CG0to5QT3GQHLG5vu3CdBJO5dHZCwb6tdWiWKvLArYAZsqwtR5xl27R5Q2N6S7Gt
pvzZdRsXDkZDOPnw7AkPzpOf14UR2ADVA9vE8nI5adIWNZ9SoMbwCpEbXqATMSwY
R+1ooz0lgITa9dMCqKUsy/a7Ol+OgqJGpcWkOIyNDF97M44m0+0evALKda/A69jg
qIcj7OXcxDleqpzolYasa/JqKVj+OYCvmlu+pdZocl39LiwVlwsEpr59Y3qHQ0l+
zlUz+TvQW93ugepbD3Y69NUtJL7MpF6ij3pyU8dOcrdJHeMHUAKYF+m2/0D6g4wR
Qx3wjP8qyBHSTDKZ5VySPlLvu+0Pu2Bfp8lbn4bcckmvOAYEpA5ivjZj5AQjZDMs
//zuaovlGoYh/4EvzgD8ZwW0t+Elyi13uYakPSx0ZKXbXLjLmXd7D9wciSEKTbCd
Q4emvMf4KhHxthmf2QlOkxlYI6vKu/P4uV28mFCjkq+QfLSnyeeabC0Vztnb4clU
z2PCFQ4jMSiTpjLvKrazrXxOz96PM8R0C64frmg0d8Bh8K2KP6kkglNBp+WUThDY
hUcYier7TfjTBVeMxj5Z8+tI6nER6XkGDXlM7eDK+L94ncd2CEWi/mf4hMRHfHNo
RNgPwfdYo/iF+v9ynPL52tZ9mOK1xUMfByXnNX5WXhXCwh+SYMcpLgrQoWwq9ZR0
L7KvwIadaTJffJZIqLwYrVpDxAF3wXU1BoHDxXHiBXt0TMQrAPLsW7UESFfFc664
vH55XDWDP9RhDK7dlsfg7Y9agU5ZL2ClZT8IXtt1YwxHY2U3+WMCr0XA+x+B1bhr
GT6qjbmMoZ6bzhzwCK8CkcC0CLUGAD723ptWzeYS2ncGB9j1GoEl4eKm2DxI7ihE
JC+SrDSDw9xj6d75mNm5c42KFbb9cL6dXbGsjNO6QYDuvEneEhEvEjvxx1GP8e77
lqyju3C5Mz1ZD8oNuNgwPYN+AG1/zw0XuhwlvwKGxb0dtXSm9ckNFf/j0BqkE7wS
PWR7dq+nSfv9VXFKMfi63qo6FQdii2yDXahFcG7ZGSLA1hjjoiSq+f2DxgVp/nTs
0x8q4/TpGCReKDgQJutIJx9dQ65tlFlNxS6ub9qN2weTsEuHvL68sl2lLA01WtC1
v/7bbT6I7VcslweKS7PRaLc1ISrqpGdYCu4IiSBnph+Yckm+CDamTNNSTLWaEXdY
2l5X9AINcPudcLJvqSC2r/ksbjXH6DIOLFoTRBJW+Z1L+DtfDwBogUxd2mLjDORZ
94agGh+k/C4klvxZLuIN6AQWVdV4V+OCpjom/08mnjvKCKiDTV9s1Hx5oH8GIJ84
gQ/QQeusKbQQ2HFgcm/DVNp/1dk0SQ7amuyGWlz2XdGD5zZtxdPLREk6+i4ssdQi
Frj4v68Eeli0YgDQq7gOyoEZHMjhqdhKRT16CGiAnXp1bpoHfiuamiaVxHRo9BD4
zHOmp1G6UEaWRpDv2mgHnFYuaKCumGf2fBH0Pxnz2Fm2REjGnjLI9QvUfRGvjIzR
IM9XZCFjI+WaGrnnPYe1kIs1K4+ERNVIcB0LpDIAbJhpbZo2W0ja4hAKtTaAFoYW
GZKQ6YTS48g0LSRocmQD1v3GhxrGxri5iWlGIn2M1o+8JWWS1RHsxKpWyDtH4Ts4
A4BvGI1UqBoyq3fAn2RuJqoT1jwBqI9mKCbpCBjsaYIIXbmgKpxpAnA5FnueGE3X
4/2YlSpvJX2OGea9+c1S1qUNMs5iOc/o9F8rPpWEHrcWu1oCPEFxc2MKlzt+AeVN
I9+qvpMsUmAghwemiFpr89UFTWWFnG9J3++14Nf4UXSFq3mlScf9zSOp3SDPYW/8
OaXO8UhSlj8f6AvsalV0aFjvpE2gJTsWf1MC027GwZKNWcq5V9a1FTXZjykMH826
IXlAm3UVp+Xql5z6ApyU299eD9wHcoB6NPPBl8P7/thYnuyUKNgXmO6feGODUnaP
PkhkgqFgtpLp0jtlLTRdrQxBpQAJxAwb+b4QZD92dJCdeR9IWTATR81MuCGjNX6H
0+O+bfR3yySX/GApKXbnu0Er4h0qlJ7OAt220xqLl8j8nwgPGMjyGZyBcvDmDO5G
2OMu/Ti3kpWgiIiZKpybS8QKl+K5nzTTMhVouUGQOlrhEWFqn1XWaKDyFYJcKOd1
3ygpsmGosazZBafz1+e4MKKa3DPSZcmoacfmGUvRijXOEgWCNNmlUMjwEUJMr95C
Mw/6biL9UC2tF4s3KgKANfPCVc4hT8Icfd1ST64ppGKBqMqJpOhAUbenwxYv/EAx
nzn14CBTP6lTn2+YOprmUeD+t+HVziiDwExkmhmoctuPEWH6F4xlEzkoG1JGWN6z
8FbEhTRZ1q9kb72zEs6p4nnG7vFf/inV9piBPgZgZ3M2n2SQMo/GfFSfdjPGyB4O
EUHFwh+uIO3Jg2hYouq0jxd55gahRh908MKIdlfO7IjqRsY0T07ma2602m4VO5nL
k0msJG4Gz+77srpnHMx+IuTpK2BHYsBtFUSFoEqncirs26nXWgJQWpZXg2tXATiK
wizk1y3VyC97709pyLXmFHG+Sxl1CLZmAwSCEoX6gzCdU6qfZPKhI7MHAuF9ee13
ZqcOjPGLhn5FL/haw1zknTsZuHs6A8L7Au2WwdRDXj0=
`protect END_PROTECTED
