`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cE8EKWNvnLuUnk0IjbpUX3na5dD4+CRsvqXbmSm9W1C8+SWPgMHxsKdB/RfBlSOQ
nsFP6MdenTpZsLpxtTAJGoQktp/GCdPc9RczULZnsdRRJy/jh6jjHjE4y9xbSWGx
sT73yYpUA9tJzTpyyf8zYpscivEGf8IEPq8ufm/hUxY7FIF9Ud9bcQJTh06xfInu
mJDv4BoKoj99MYVv56dZU3Za9V1uTGPc7c5aAo/bqeVq/iyoB6occazSIRcXTZ0g
KzSQgG7sLLhMqHvPhB7ktmfzCnylSEpFRduE5sFLvCnlhE7D4Uj2QJ5/OyL8Hx0l
+N8HrqwiKsjILjXQz+lF9CuIYcMpj3OOA4mRAdjMBCXvJGDLydF+ICPT9R9u+uAR
jJVAQjRtzMUTBJMDZ9c3f9xWhG3BXJieaoMc6mBQ8wHGyaI+gniI1ayfN244AzEa
s/yJSuDyN9EGW/CSFQ5EVhOBtx5+sJx9pYszTI135KlOclOxT9AE1vdUE1vnqKqd
mdf9aJv41w3z7P64n5c64yQkEBewOQn61blSgf2UZbIjkaLuetAu/UJEPGa4+Dkf
DBhNgBQMIxdf823oIwhmfq/wkcZmiicNwt6tSNgKXQ5LCXq9eqmTcwArX046nN76
/JkCe7NbffWq8h0a1jP6b2OGiVv23HNFMwv5tZM+i/HKMs+Vq5ISOqcNjfur2vZN
a+qy3Z0a7BNWtVGBDgFHBIJQGRUUDAI6ghJp46z0A8nMQGAFAuvblQjP9uhSGJaB
r5o71Cxy7sQjmuWYaZgFMQ0HX2Boko/GL9b7Ex5qKTodHJBzyhKt6McpILvpGkh5
bAneEPAS5QKT7HgjPNkFlA==
`protect END_PROTECTED
