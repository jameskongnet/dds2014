`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CuMGA4AuzClcS8wDRci22RhrBtDhLE5BXBZ+oDJ0cjiRMv7eWWMIAZtCEfyKH+ak
5v9eqkDPen0oVBvD7Ppq/A3vyY08fukicwjdl1FwOxpVV6aet+3GAkzkMDYNTR3g
s2O16u5V6WEbx57NzvrsX0tU3x1wZxrtEE82BRxgM6uUik2Ap+E5Nx82ufcdEnN0
TTXH8yE89en5LEgf1r5t37yKlj+96r/StoQBSYKFYaPOZDtd+o+kUTlOLWr2Gm+H
aNK44Ach7aUj8Jaa96DaZTXhEWG8Ujvv2g5ktW6Os6p1U1nwCoaDZ4LK5SyLAoDK
jZGd2DOTshDTXpXqLYQLRa7WUYPHIgEYcUB4IlNjwkvQwVHhhkjXQ/6QBkvosd9c
uEsO4/e0BZoHVXrIcCm47KOSsGB389kGPLWiJfcRBXCHm4KsaC/MbYvai169hc+z
Xwwf1mfss3M/dtOHwUgqyTjkahzWsvokQsZj+XVqCCtdOOk71P8acQuyc/wXcJsO
d24UyQm24IHXYtROL23+n0xx8PftFR6gzROJ/0XI9KqO83I1zUucoxVkZqvWEhPc
ab0GRgsvUDk+esNg0OFUb6pXWxrtllcF3ZRlfYkVHvNzLGJjwDoDDfWhOGdMsFzE
eho2tAQZMynzIDPFBIu/Nefi07MMm3EWIySdT1AVRj6a6jzUj4dM06dtTQQ/wpL/
tkLOa2lJQ93UNPiC3ZKkQigUXZzeGriD9gQRXpyx19AnnnvqmL7wdr+vcqKTcan8
dZw4h5aRCoAB5Lkaih5Dog0v9am5y1npj13XC95uAvauO7IH+8CY3oj7G0w9m9/h
pqSgWP9FWuUPN5x6jAvqHeGQSGgfaeR8zSmCE4JC2PUzrVnJZWK7ZCDoZ/eJszWG
owhhMPFMKtnY61B0qKyfdU5HPgkGwBtC0NojPujvHDw12kz/193C7g6FseXrpxvb
HMlju3r10eemN1YmkHoEjwLUDYP+ezFtJtW7VaO0jz29C5Rse9A1ba0LfMlURCKf
P0iIdlyLgyBT17JXa6gaTEo76ME6pkpWfEv+spLRgKOKWwhUQqvRi7s8bQsmRbow
y+ysG506IzRGm2c5yPAqAqGnOamlFme1+EbVrH0o7yt3jCbpydjy7jIHLQFuV0lI
nhgTeIYUVMXlFmGBuRKtu2R23hnvBBlymp0mhP8ZwNj1czuCvMrJT29jsioWvAA9
KfVpzKfj5rhUVITIpc5DPeH6iIrtx7o48bnH5UEuo/iahS55YzDqarGN4GXI5UTq
V3IDGDgdLciVfRadhqk3l0c4SRwZx25/a8PBl9u8v8Pvf1DvvuiwDBMdm/G40Lah
X/gpeVAmBS8HIkW8y08wErEG/qiimuX09wDlUFTp9kLa2Ke99LM5YiuqOb6XtfeC
3FFMmEBi40iyi9Zj5BGawePiOn8rjePamIySZXIBZRF9lVAvLxWL3G8wisFM0Jg7
t509RtDPvj+lxAeak3BAPeJZ86mwzHnIWqiEs2BF+DlWx0IAn5+4u3e78jI9F6j0
x3kQ/HQCe9wm3+ZU9FW/DX3K/sY4bLmtmz2JpdblSi/6rn3HSLP0Da6++1I7az03
K/+ksVoFhdYUldC8ct2tKSLnN1+VXnQhNiEa9/uH5oH1zZ/fh4vNyq4aAHO/e0xI
aZk0phPGbw78dihM+IuNH/8w7DfsBbXlCkGEwH6Quz5O3sEkEl2/4hVUNipAzbRy
mH8nNhFNTCh8U1DzZCleTyyFnVJ/KEVYn9cZGMyUrnvf8+y9ko/8HJ5HTg7hGHfN
PFv6PRFOYR1YOVHIhb5oJps+x2pBMJkbbDLEL8FMd05I8t+wJbl9j/ouYkhzQr2J
WydYnRjJ7P88eUCHFEeq3YBEQzTUJELC6YHbHDfgKGBgDCg8DRVShJ/y/axm/0EZ
edRJC/eY6i0l4zQlgucgXlTgy5W9g1eYA0LE96mp9lYYIpeyjNTgAiUMfVQfSCV6
YEHfNkmPTYNI+irVhSffpNlOOcuM/EocV6z3mqn3Y5IctkThA11bhhmjo+Mwgiwt
Vvgs8l0N9pXTD8U2Gw+C/a9EWnr5OkCTs2oAVl3mrTVEjp/RXOcrT+Bc2jeKriEJ
MsSo4OcVcyQkHWO4R8emwSnFZ0BdbZ8of1TFN4Gvj0DqZtAwR0EboyZgTs1CFPkr
wTQdIu8G/F5cmJ9LYsCVNIKFcoTQX/9J4iGIEE3kr8SMV5Ld7fbxeS8aP6Vlz1uz
uDwApbcWJuS2BzWjB/nzSS6K7ti+Wy8gyKi3ClNfGls4V6cFuZUGj/znhK4/8QdE
e0a2NkhRwt0ddPIS+/qIDvMVKzEuin8FWy/c7HMUp+xDA4yiCLf3rQ/VRpTXe99q
rCNKgKMukALOpad8dXXiRllrSALS2+wMMPySIhqwsL4t93L0Qw8HjR8dT5Qt4j/V
j5xd/jFFDCuXOdnZhp/gZ6ZYAFzmIYWob+yPpIVikPNPLXF5IJhIedRcoXeOsVZv
ayqmmWASGzqYBuxjenCLLVep5MGSOGAtZpFEbASNAsGtzJEgt3UOhLSexxc7Ili/
EllU0Fyi7KUgGFYzcrybR4bdqntjzhOw3dXxe2lQ/gBuQg5s9+lmoxfzOKm5uwRr
hBJf5QVf7V7Zi+RXS0uwQ7f03pOuln+fnChQZEwR9LTCe+fDUjpvv+u9IuvJOAYj
jTHsOG2SOcNix6uRFwolGFbxfrtUWuciT1iHYkdv+Y8qlg+69sIp/cUJ9myttU3i
AS5NbGjGC7TcpaXfJy7s/WvkAPleppNAVXv42G1518otokVU52h5yfUqqpdj672O
G4X/KwdT1QdNNUDhZyyT6IZNllD6sbBJRDEHy5AdQ9ybV0sONRFawVSt95apJZ51
aezfOb3/I2SKgvjbV2+LdkbssUxi1l1i037GmwTxvOxClQJX0pHrqK0ZPEkTgJFb
CwP4CpanfBxM0jtsbMMqGL7S4Z1fjFOFWRTBU2IjGBjwN0VQssi7IqD5uzqFxfdN
6B0flAOYFsp79mw2Kb+9+/in606Y64Ooo9Os/ejQ01YHjn5RmfSqaF4Qiw7heiAF
XmrPeFB+O4w90STNiPFpf+6iEhCkGblXPUHqaNogi9vkAEwB6e2ZHdF6rYnrwJYl
si5CdlQ+O7Ozv4B4ExjHpd+gBh44BkbJGYvJykVfVxhtqlbMLGB8RqrcNOjWPbih
MV7xGyIVEhoH13DtsR0fAnLoHcKDxaQtGM+bBjojj8y+wrQv9ZuDBTpTfPDY0HU7
QVio6/wP5ffSr54+0nEN+mG+0UnhD4DWIw8Ft3bTvYGUV6M8RV8X5lakwBCUjbeS
qhC9zEKX4jm6lsuPpW23wVfucl3BYd8lPXlZG7hTnNe+oP/BFN7lUyG+r+wPW8lo
OVCof7TgcNJjdvXskVprijy4eDpSSmnhihaPWA07RAQlpQP1sq6cfIZcEU6G9VHh
KNJ5bGQrWEAFOMFNHY56Cq0J2abdQyri9Mx5WR00SlHDEhekupKbpxQGzP7nA63b
6KaLthJt2HQIg2K2o7wbKlZyDOiOdJMGTNO2slX8C4dQ/SnMLBlWzsQeSMJ2mA7U
/8J6lHG1vwozQQhDD8EchZlzqdTocQLBRKiytekO+o86ahBQs1G3om8i6OtMZfE3
w3biuiW5Yte4MUVWP4eMdmWkXjge1n0kH8SnF8TzQ7kgXSh1BHHCm6Z3lcGJbgjk
v9X3qokyxiS3fNMnc11UF4eItTQT6Up8hNuO3bDPMsnM49MJ2RbyKWbboG0sUEAg
kpiQjlBUgoFbL9WQXgcwT1gSNzo0mJWgrFxCiyEPc0N+SiB+bWG7AXhC2mGfiWdZ
H01oCLjrB8prBvwxT0TEsz9+M7oAEF258qiEc0PDqbb+n+L2powG2qtRchJ3HBJ1
QOOj8CGaImT0lmiWhgyYDoLi9ZkF3zq+5EfveqTOWU7cF9wV3gYOzffgoiVrWBV2
EFN4lHBc2iXC0ILtHQqmWA==
`protect END_PROTECTED
