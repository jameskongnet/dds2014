`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJW0EFgtnQPvfvXR7mBYIOH2j4/SmQp3EKb8H4B2dljQ/k0rRY92B+dLdNPDE7hj
HxCBGs4l8tx1zrv3HapnquAmP29SjFW4nAphJEZWOyzbUvfyL/ehbpdHZYH3xE3g
dFdJTPkSWl3YzjpqrfUCVkObEzKbQBbDN1xUepZ208Cza9AEotV4ybHciQDexMfi
SQ/5E/pZ5YhEs5p961hujlIasQihFv6p8CtwBZkjh66lNTUsfE63/QQ9UEKfedye
T+ZPHUaWV5Hr89R+ce7OWNSGvS6lfViq4qFR0V+t0Yis/6xojKd/MjR7ESEdoOuo
iRFbu6/LW5kxyxvGw1H1dKszwTeJe4ObBrWBbkiglG3iw8LxA5SMgLfH/1H8omoB
khxjCm+WzR8P/A/tqbb5hEWmqUU4YaKSGticCGmfv9l2u/5tR6ZIRY0h7A8AaDGK
84ULx2Pr0sPVb91QfnwVc1U3gaEQ2ppCdsefzy06qXzqD1v0dri5EpZAZERkfu2d
OoYQGhuMJLNXsCkV5RNyqHnplp36b8D7o6yUqv6swFRHv/EZ3CoX3Y+/ww+WTNHm
yok6pvOlXU6ORpFXWIMb7MU+fJ3cU+LZM4RIfy+kVN6jNBO2GF+OiLOo8dun4Au5
Tns9mKCbixHlPuEFO2ybxJA5l0HYrmnc3lIuyg3aqurgSoTedR5Zfm+db1s14Uur
jz1GsM9VlF93NSdyQ3JWXQ+LRXGeODbDi1o0tZAnJ7s4MbSjRP3NM4r5cTY78tsl
eg0tSZNfIabyn4oPgbu8nD5yyWwxNG1S4IwZhDTOptprM4q7ndS5MzLHgDz/TmQ8
TZDxdpLrXeZf9rdjCLe4M6O22hCWhnQ9pN+F594m4wJ3zTsyymeFkl5sF0CD4OQJ
gvgjVxOp5PmEFmK7hrUpECkaTv3G5ns0hxULDHKaOf7LOfKwK6MdRMV2//uSLdRg
0g7IINuArG4SswdqzfJKFb1XAuVd7QcV07FdUMi60DGx4tznKspgAO7xuvx6/I/H
bCIUlCxf28SEy4gudLYRz9Hk3cKLzp9UysXW/r6EMIMyVXtWTnn9qFlOQWZ5lY4f
N7kKQs0/UjvNJo+KXrwcm7J9hoo0fcdDvEPSd7AzIL0YR4KskH+hKb80zPrV5T0q
4IJBirHGaAJSrsGicUh9q/T3q19aH8chhvMGvwB/oAJAezoPcuwgNz0YIjCRnbce
db+vLHofzr5tdD1H51URL/hLUp9nIFErD6eCWv5lKAUzr5SeqdCrFaa55c7EdavG
sLv0fwNO78Sx1vt/T7NHd0HCIMGsedxhSLCcP0fEhGc/esDs1ZYDKuhr2Kj9pnKU
lQkNmSg7KYFfkMIIkPieVVwmfaCEV7hreCzAFscZGPTftKMxppd6z4RPPLrwcjDA
0mKMWg0U3xfeBNDKbjJ2i4Okgt5Jux0rt5PKa/jWpIlEqUtXeZpeP5b0B6fnrEu8
XMQJoUtanY7zRLvjo6jnMwxlH15Hz99FiDW3gLwC6dNtOTC8ALnDX0q7B2q+wyyt
6vrr6Vr0a7DpzelBINDwninK5xz9OGr8pDBcvOes526LADEoQjY/Z9seUoUSID1u
QBZgy2mf1f5/LP3+q+IWRzngcIUVEDaeWsNL6vFj5u72byQfuNPJMEmYynreWdHi
3BfHoC+iDpPijvWvW0Cy76wncF92QqFuaCmW/NTMmOqYECIXiV++GkgQM8+lHk9b
kpMgp5aOlvuc72VTEqIUP57KDSIxaEYktCI4jvSgLEX+b9nVcEoR9HXNAuJLutXE
00WxpZOrlJlI0RfTGnfOGSJtWDOWatYFFrLZD7XEWpUJpesr3GUhwzYgjjTpnG5L
6spDAvXZxu2JOFjgYOkaJoWizGn0Oh+9oSc7lumeODeKXzC/SItkGFUKWkFu3Wkq
AzCuG5GgrJufp79SFLZnXWrmW79XutNTM5ePvx28VPej8nsFN1GPrcMzQL3OtQMd
J2NLa23iPX9BkAHLWeMFrCFtsqy6BFaWPasmyJW3f9uR6Nrw0em6mz44eRXGpSho
Zs9c88gAEdTud4N9Le3NYVhqWfwHjJq1QxfzilHyFiWHCXcA8sXC2XideVxogL0o
ZsuFjJhjxwNE3Kkjjnemu/X5Vy3nRUggifJJHL4wnGDRpVLtO1cU73SBOamrYDue
3PNO+M7WyGUaFZaAeN3+5Ym4bEt0OVmnjM7NqiOXAVQa6GmNhH0uN/XJM/yTv7Rz
ptFUOzvuv2ygTTvNs6N0lJoajUZkqEHpe3MDQANSovp317qeTTxXVHMrxmvBelIC
xZ3tXbMv9IGG1G+TYJxdI4+HMw6O7h1gZypO/17q7ulEv2ooooOHCPOlGNAtu/pJ
NiyHm6UKP4cplbiH52+PonyNc0LB4u/nnLkBQx/Mw06e4MTg3FD+C26U1a1x1hFR
9pt3hYFgUavjvlkoyimyfQGLyRrSGauWt29pec+SPvFOQGUBpMEyTaPSmjvEOA34
zplJxoLM6RFJEXyXB61VGLjAmPTu586S0T8afVl1AZtlFBUOWni2eYgM7ictIBvj
DXYbqrH//mzCT4HtP2ZT/MPRSlVD9Q5NM65JLveqG6OCko7597CQNqbgWxpKyyaw
9qGQu0npjXuY5yRrUkIefGQ1oUA2mj68MlO7JNKsVfpyiGDbI/7GDzKj49GNmmip
Y+D95R/k+YlN79/y+7/gfDAv6pdSmIlqvEMVMtmDM2SAl+GgJLbaQtG7UvrWJEmA
eGGLjMgjhNnwXvNkXTPeLxLGK0+ZNXZ4VbTQYCDsN/i544Q/NutqlqYqiuy3yp36
zSUXibNn9A26kfvp+ltBnqQ4l9yJft5r1W9tIWJEx/dnPbuokMH1qAXtzcNhVas4
QcqIygaBs8Uue6C0hLYL6ziuOPJb6T139kdP5kj9IYaJUsGqpoCH+IKwPR/lOeVO
nl48P4rqY4q0z5Bp0zvhQ/MkCoy+WURKE1alnVGmNqI=
`protect END_PROTECTED
