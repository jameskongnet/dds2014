`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QNxWw92vRqnuBmoXoDUpBAD8mAbQfDjDMUtje+mQzOWiLRvUjqrUcbaDc/3xO1CG
RZgRPiMLHGcQ2EKrn4WKrn5/Wq1JkBA1at3fC+W9zJ68G5Fbp1daVnlVw58h/UtP
30zoRVWvzP2ohghyYR7sLnkVRdNA1ZaCiKTPqGf3QrE6RiXsXXXA6OkwIfHg5lm7
KVhcoj9cU0o7OUqClf/kTzD/PM/Di6la+8cK1606VjiAj4bsA4dtyK3smDRGol6T
dRNJD8742tKEKu67VPkq+lx6DUD4rbf9ZRuHXV++VLNcaQD1lqJKq6qXCU8uOxyy
yVVoboBiEXtnG3avQX/ZDhsXRk/BMy+VDvFaCdXKmGD/pueys1dibV9ieAjxuD5D
2GNsokio00ZqVLkzTcKjzPhO4BhBv0JpfkPuwTT5sugVOAQTBrmk4VOG9Hvokdsf
K4C7ic6XQovl719UQ++pYzfJNDiLTdh5lNKvlPYT34RTRuyjFPjnRaXYbuynHKLB
RdSh+uEsCdroZF+EXBI9fMG7o1gkwvFdzwDY8NT1dKEOULJLrpWDdlkdzG2G5pak
94xUmFMgb8KjbaYHcsQL75NSCAaLTDdB7BkfgX92SGUhJl1hQ0f3y/KcKxt9wlxM
e6sD5Klsq0UVRD1N4/PkF7ZL7IAHiZs26Ze8iHqZhVxB/W/Smts6XzRN395dEUm8
aljdR9SkDxBXCxJ+CPkr15YN9IRCDDr1D6MnCGcPDe2jwpQhckpboumyR3iekyKh
XXt3Didv2g2V4MOp8lDCK+09vJQX/AjBymAvaPczwFMW2D7VoPlyNepTqUAMZBlK
272hKZGdbkYg6JX6ahVioIOvB9kvLszOe/Pdu4jGGQ+TWp8z5v5ERmvhRY6R/BjP
nQg0Jjd0K+kK9hoVEC6ebiSFQCWvwEBchvGptm0/qnC927VYdt5qrOVeZIU/sV1z
PJUU1HNRD3Fiounwg4Z2ez/VOaTLlocjvJdbums3/pnnXa/qv45fhpefGI+NBbyi
F0VHD4Z/JTgHSBB4kGpHGLBlY4qrzOb1er67ou+81nqYhOTdzS1w4YgxMQixhZqU
y6r5U7AGsixg2Thn/f7WFekoe/nyz/x+d3SrRg5inaOtRbAu3RhqgwRs6iXfaemE
fbQFbDrqi5VfpZufhNQiszwwO2ExO2bCw9vCpeG0iNCimVmNdMfjsDbQ5QblK3e3
jRv8di80YiRpGqjHPB/LEvolSKz1R3/U/NlsRvZMrLpllvCRbUAShmNDuXvzbGiU
39JSsqpQosCacJNJBjzC4JYe8MDUVb9A7+fJGBSrel8jAA3F1w5FPQXsH5dl8xOX
l7nfbJdokmw6b6Y2PaWzntGT72cD4gQEWDda/osI6bbCydUbyqgy2PxKY30w3krM
GCiFf0tOU/w0V1osf0mEg5lKAq9+Gjuwcm06rET1vB/ZMbcmUM1MeDv+e+sUpyWv
2BimcNP8ndFekp74gl4dRSHVs9eZ3ntZb2V8y7iWM4jy8byi/n26bdHmLXvICyKJ
++0HHdE5zHO7vgH1X/JUNowuBQJG4N0eg1m7ltFzO7Yqar6xvrSAAko0fzap1eap
THOh1eO2YwQFbc9avoa1cs8Cu/bvdHly/9OgBmgL9tUi6/sbPndY270ZqT3bwacE
ufsGakZKo8888hiDDjL6VjOvYZiotgFGXsczI4O1FHq7yROQ4xuynzC7kUEkKANK
hQ1yxLRVJ1d7mVwv3xVTCvK2ScPKAGIfrsAMipvBEUenWaJOAdQ6xqwm5IO+NUDi
REyn18HFw7vVa4bfCFaBUa33DIEhDh4T/pbIZhQtAw5uLbsGsN+tFW/fc5cWEfbZ
jo5+R+GvIgOjoMAUfwlussrNmGwqKqbLTnQIBQsIQou9B8OYzAbnq0BoskE6D2wS
OZouGnET7hpRohbQQw+va784e/QKkBX3D9G5asq9vnKLQM08K9gQEElfNrCD8Bh9
j2qxRsvMxKooKxVSyQgEMWu94c26eOp93UAwk+wB6DPqqwlyRwK3tL2AA5nE9VlV
wwLw9jCrwz+Rk0kCmwfeV3jtAhXzV46+BQZbsYMqQkqXDS9OWx/w6iAZ1cVQ9k0I
6/iD0UdgDfVBhtx7oDVkgbbbHVgOo7VkZ0TTN0ifNu5oPHUuEAEn3eWFgvxVzkuU
UYIBxM6P0H/vPkqqjPUaG73/RRG1ksW3ndn2RX9VtnNcVfIxvgkSD34NE1gXDZTQ
XoNTizGjsSlfEUWyFbGYSClAWJNosEMRv7iy20JGAShyibe2kxvr9xidDNuvt/ih
wfpGRUTz0MFcyMaB/qNr+mBUTH/KTMcrqZH4OkoHJlWNw/4sx6aNavk9KxagC4He
iX+0plEmVfp5eVl1JGXPYIR1+5mvLP4DDFHEfPfotXr5HE2eJbIoK9Zhuv1zuXwB
Odj92d6icYEdZZ4Zw2E7DJz8a0jPYIuzKQwDhI+Yb5HKa2F0VdpMmAFmzZooJ+qj
Dg/Nm8NcDaHle2Px7V3Gcqc1TIHPK40fKPrpmzokCk+5REzksjvOtkw9OhkpMdNh
EQG7BMcT+sW1h8HP08a9zTHiToNTcJLOAGUMRqA/R0RVOTuL1B+2zPHIxE82grAP
RR7tDUXEcoDCn4bLhzbV0qvkIw6KxtVrpr2OuiYNYx3SFpgkqA5x+QNIQ76vnp4G
i0+O1sGaiNC0iEyVefdRraPcJD207LMtQuUSV88gdh2PtaZVjMZi7LblZu3Zycud
swLptXbSd9A/ot3sdBF4JabZJpsVt5vjFauyyh5h8GF/8pNJtZwe6i19qOOsodt2
8qJ5KLtmnRglHPIFKBs38678P0jF6tn+T4fqRVstkvEv4YWnocKBxL8vYsIEtBrA
f3FxLkVUpiAxSIbK/V89XTZpldeJleRnPbzZNK+/+qbzpGqAX3ffQ8in2ncjNlA+
0ICAkBQh3SgxIfs0braN8ySCKDrILp/wD4kgOo3AIWIyTydK5ygc3PYBGFUXZ6ma
6LTAlAC2oKCNAn3wX6GtXzEp0LiosVUt4ssiCYhz2OdonMFG2SPU6M1tbI3lYx9x
RPGjbYwiQ+TA61WMToW84I9PLC5SJGnDtom332FxLNfWJhsDfOJy9k8OF9gT348b
0dprEIpaQ71urZmRitGxbI+eqx73GYe6G7oTpGr1uEHCu/ADHTBzRjazuLnQMVLB
peZB7aA3dc6VdHQxSulpZ0UVCBtm4t8TyKLu1Lxk5Sh3KL0YS8f6ic4s83Ojrh7+
tG0WaYxSMlDc3qHBz8vuqrLm7iTFNpOmL3kNbzsiuU/VLtJecbE+WWNPCoVZ7VhY
e4pJk7ITPPciOTKgM1DFb14AW7UxtL/Kz6LInc1rKwS4lWMiNxkvsxhP7VBfAAk3
yV12ITDlKD4viU0h5X8smKyYpht3B22vQFMpEUCi+Qc9orYA0pCkUuLsnPjSj4nY
W4NuvNE7iNpOjRyLZfmKUc8zlCq3t+XmWifWklKVT2JuvBsRf540JNYo+Aa9bF7g
xtC8zeryIxGyrl6XwYzrlsX38OW598KZdCYMwwsb73FsTuNAbZIf9g15Gb8NFeip
LrDbLzemRK5XmTXWfRAjWNdRHS26OUaru54jIIuvMctRURBspRaJWnUJIN8YQM2I
ZAz7hi4d1KAks5W7hhMOWYaG6diGJJVclOSUyA9Fie7Htc7MN6jesaKQCljdxIZ+
41VP6QbTCPpshmgdNuCQjdzOvO8HPIFSrxEYQLWvSfwJ1f1MUtpeMtxgTIWuWUUl
G5um40bc6zPjG12GUof5KGvXfCHmOdmZscUCdvJwPS6MlPSEarmuSeoVFZRu2rVi
qDadKLjfiXAILQwFmNrm48qjG3HWdZz+3rUgESp/5C2ycD4TQK9kbNcalEfw7vmA
Ey0Xk+DukUtAQ20WWsy+tkOvOfnaK24IhaP4/tvwdb6VALlWTfYuF0i/tsJfxS3v
JxuyJwQcspyP5rLPXzG8XXq/IuCJ87XyKhq2807OoFgadMegQPmiNmkBlr800dhm
FMSXvtbFhMD+EYHH9WW9JkbZ1LR49j9VjyWPSemlNPLQ9fyvutcYhNDavwfzqt0Y
ZVOvJFhPJgwPovm2AtuCF950zfAd0i+OwBOSyJkzx7UCdwp2fZ7mCexFwSIqTMSJ
elEKAuGWg8cqhym4wz9ByKEn4s5hQ3t560ThboRl+280Pxis/iPEq44QiJRShd+5
mzUj/ndVKBdtW2RdFy0wi+ZnZEfTnnU0Jo077sR9vk5hfrh+zLgop2Nv5UXu29Ng
WgIJEWYa0PjHBLNukxCuAiYEHJb9Xd61LwA5fc+DLSNz4gBw96UnS+HHlmI5KYDt
e9RI5LnlTK+HA1QG8mUKqWB44vuddMd4k8IlcpTjhbNPZb2RssOTucFh8AizxT8Y
3M52ZwcyDFKwBScwfFqvaNtvdGyQS/F+3xTT6Di6lbMvaiHREafJ1hNo0IPc0L3q
x8Uy4lqOmcIfsVvSJnj6PL+jAmyXiLNy6pN5wLPpB+f96DkfZr2dvKMr8pVYl3Ut
/s+WYkfaYWKqOZ+haBLYADqaQWPpOa8AIUztQyOhmQAaOsfeCtCLkdiD8kiGHhHi
wmnUQeBRUbrmYf9f2ew4WHd0b2hC0ll/txD5C8gT1GFzaVhP3z2/JH9ZfdpbMGmN
RK840Klw1Q92+hLeeIsDU9JMbVY8NP/sSQLB6U/JyoPfiMa0UHDe1Vpp59JZAks9
TcGfuET8FZVRCYcDYXCx02hieBGJcfP/XoBZr6Y5lFWJ2VRpaCNhjU8ULO6yATQi
ykV/OiO64sq2WMt/gtTG93YAoETaTRksQyjPRgtogWD60NgQa7/gBIvtU8lNjhec
rP0drCHQHUaaLuPJUUZRs+VIHiJZ0pSN29hxwG4JuBtuhmnSIUTivAY28Fe6tO4W
QgKsUhiaGUcU/XdRIm+YSMgqb7uxOgD0DObFJiHwzAjf/Y3PNNR9ar/xvHn03GYw
Yq6+VqhcOBLSMx0leL0STnKcAHBP+E5YmOe0rN7nR+wXnMwGIP5cZMvMM1bWRBGm
wi6iJfMH2M5pln/mjppEPa8jpIseCN+X7nwMDpQLjr2urjU1vr0Um0pEeTHZOyLf
L23LFIzopC2WxSegmt8QzYVQ3ZhVV6XCPJL1CcqLyy5P+aK8SEdW8f5jkJ4wXk8G
TRyWpk8b/nj+dygTany3kVlr52Vpm6Oc2apgsaMSHG/TWNvKcFsPXfNKqVoFb1Jz
xJJCfOZJI9vQ1FOrzhvKALE2KDlyRrP+xBn6PrbEUmyjpYC8hzVt44La89NQfWR9
AfFjPhxkjXBzdX61mB+o0b2ivdb36TgssMVSkiGvOtHjcaIfvsoifaejSKv1vYCd
KxHnThK5ozbqreaSApSCByWXy0nJuJ1rYhplB66dE8km5bNo8FzSSSrgcEm826o/
lq7dFkQS+eD0yuIZRwakweKizDjmf66owH7Ja4n00k8irga4xezv6AskPzYoAZ4e
gY+YP4gbJrvIYAYiIwfwOWVlUBh9hkqE0NuGV9kQGJ08g9WmX0cRPgALcZcWh1Qi
0fb5VYwURfrB9tdM3wvkwzHPgTbfpawe4n991/j9t8RMWKwTKAdCdTjVOBv4/360
e60589hncfOjcWdxkhhIvoCGcAXpRaxliWq4zOJTZ84lS2H7baxeK+dJN3ZYGJXN
XtYciMOJSr9EN/D5A5BtlG2nrON460jvZsPww0WHgr9Xi1xNs6tUdEJSnzkAkQIa
cMY//FPe5KqUnUew0KEbSltlk1JlB5euuRB87F6xrsSs+18pDCpgG9vWi5NtXVZM
KO0kcgesO6+GIpdXNBQN/7In4En2JuBYrij2c3F9VcqQHU7/GE3SlL4NK0riHgG6
oPT5viEUhg5u3KmnopEHjPXE47cAwQGBI5PzlyDiWbjSwzVJvcauDf3cI1GL2SG8
lVRzEZFDAMb/yCj9QcKOgQNK3BSfsrFtUgnWo3eknTPt45EIs61v8DamzhJ6taRQ
wcXQFjLecRs3MrSJKPI5OmPEIGA9vBwqJDERTwAsKjYsLtyxhHmVXDfLrOawpPQd
Tb76MWO9bzBQieQ3AwEioIgA6hzDgl3uz8ACHm5pOhXTi65tMPz68SSlaKGiJUMv
CCp7YpZAz3/QnT706K2zANPFUZwTY4Pgoogv7XywixIg/n331geOqPQBbWgqZ2b2
Y7zB9lvb4i2Pq/89+F07wv+AliaH+F6xsJ5z0nLcJduDZRh5HUXNwxCsVAo9GNQu
Tsxntq7aXsvH0QsGdUTG644KXqEmyVyHyqY1YH5EE58iRWT1HLjBo3cMbHgLm0/S
0zfti5GhIPqJp1zPAVTKH290m9onc26GFmuO0p8IZeXQ0rDuJRIEFguLNpqlDJ5S
HQuM6ZrfpPR1ldNCuboTi6lCFpz7VlMqVuhSvtsAzGKhcC0YXyRWhyq3Z+tt2435
Hy/I9nkdidpZbyaLidZhn+Bkou6W/BrywmCcRO3d6aVqv4ojQUfnUn5pzU1xGs5H
1FR13oQcDrKhYZ8snl+gxEvldimrl2IDY358Qi0jrzbMP3w0whAcQWDj31TfeDSP
hB8uq6cKJme7f1U7gBTEuIElbGPyVr4H7XW4v6+HzFk0+QZPCnYPkhTc/A4CQ6v1
qVu5ZJN2qBYY+T63U3ciWC5HaSSKJoayVx46LvCE+zwdmK6mL73e5YOWxCL6RpYu
yK2ASmT5r8Wyv7zRL4eeU9CLiUnEAzAhGXEMplZb/QEypCmJitVdQCxvZjbsLI3b
C62D55osxWX1YQlXVjZAZ/7OWThIxJpQpK4OCDoWb4+dq6dfwLmYyN5eDOOkwvXI
2jwBWbsHoJZNXOBbbDiRSkc4Du6wta6QKJWUVsbLdWNUTh7JviDlDFV9OSfkpz2V
JNUJJer25Y0v3Ff8IZlceizNn0jBTB9tUdl1zif8bROueb8YCurgC3InHj4xEo1j
Q1/tDo4BdxEvPVLgd0+DXUjzOECwB/XAjS6WOhKg/dHBQQ7ghLd15g+WXckcM+KJ
sGYSHJ5jTvssPF4eslOApOLz9ZU25jlsrxeMtlrTJY5ZXApy2EVoIk3zDJSCa8ec
AfP12gJXxFtfv2zKK/85YMD1ahj7MX1ufoMw7wvjS4RIW9l8PbMsaFbYpEPEkVNu
KdBpuN1l7MM3vi2FF9MjSwj8pcTQatTsuZsr+6evc1l97W2UV8rcJlLlUJ9KyXb1
xsbau4IgHMHc1zpf0ObTdbVYY24DPEMQLgW340tg9PLeShTQQhKUkr6ZNgoNhm89
BCxawtH5MYxju4PbntbeSI/nuX+0TEwhiigfQ+7DSE16nzBPWUlarmOTHXo9EX0h
vx1JIUwOk9IaxnMiotryvDK1EE5EpUVgsx8dU20u3fH03qnbGPOZck8/IMoaRTNk
ve1Y5eFZstpaqvVxnq9L2lwaU+Jltq0yv8HW9JCHy5nDqXwJZgbUkykw797Vnsjs
fX+5V9gA7D59BvAVR0BWMTRdO0yOmmHovCoYVo5RWBy+qYQ4lv5Zb56OIknQk39G
6JTZOsW4Uq//ZDTQ5Jb2dt5dpaV9+bSPCUPdSi+s30wxHVaovBrT58QlyC86lVzU
7YbrhMTMna0O/IqasxDDlhSadH1KmrnBw+TY0dJpYxZAAcUYJW1DIeL3NnYaW6ks
2UkIvzvmOsLE2NC/9cc2fJiuMiomVpm6zVddBNe1j1tddHhXuoJc1kDvPgITEU2z
9WEv607FFEXlglkA4TawPBOS43zTcbK6LVfRXshNtewzR4IquiEbx+ZRVRwUAlPp
RyHcG+zG0rqHcuMB5OI2kDIdaoH6apbgO4eb4epWDhLT8w4DiQ008IxCYvM3QeOR
TcQo343ygf761g1ufdnEJoI0aAkdNKqGLDyU5ENw8fwTV6M1xV2HUglLJM+N2tTL
6yjPIWKIKD4k2ucohFKUu8aia/OIOdlXkdUawxuEMSeGeTIkyIV8vNpV9PiJEnY/
oBDw0A48IJkrdo0IXuKtvrwtPsrgBuKoe8YL9V222YghTKWLOWdxFBWl+9fOfILM
LTrgvCbNl+qNDSOtRhq+dJpKUcwt7hX8hyd4afI3M1OFEtNgIi5XM5TjZpTmPvdW
aZe2EZYWPvpksnbIVABmK+qRoM+6wJz3wd9pJ6S5Ev8gRhr7o4XMEae179V97xSC
cySO6fDVaGq8E2mjGhpK8R1/BnhIAjikV8Qh6b/WxlzrGyi31b4TuUraUzKelF6Z
Z7PPTaUo6naLQQ494TRHExvrHubqkXbTQBg8dShw+sc8NCtz7tmie83ZbPtxfGre
MK7DHnAecMWYwIoEJcgKu9kBCEVCIN9qIzI/VMqZjZ14cd0cM1LtXq4a0byT+9oa
4gc/dgSDYnI5GQpQ4g3+J9n/uZs0mSrZs1OP///z0p+2VJ6uvfQnEHYuhjz/bHw0
ersT8YOCboaENtpayFYSRLg2Dzv3b8FgJ7FnOYu3OuGlhHEiqj0iOEXT9wjPNF/P
IZEt02u1l/KJUILsN8GhScLBJuZFAzZ+gc2enS/gFRXf108Z/e9ryvHDln2BkvHP
HuQY4AcOtjNXtxwZjKl4XNjeuztiWBRT7bntmvOuNw5U/RfLHel3QEN4xBgTJG0U
qlbTmbjczpX+vn6pfYMPgkB3tGxbf7SVl+Bs4Xzc+iJ0lD9IwPTIhmhwDCET9nBm
GwaTOpd1H90Oc2uR9632X4EOydFvgQ+1svRn6LCdUWgdaCpsWWpeSssV44SuWwZa
jWkPcjODXQFD/ZjLNNIdNx9NAaM2vmkw2I+FLu2PMY6h5AR2/dHmhwjybR/8379p
ZM2lnwKttq8cnNeDzGMRNEp76ziNvhzk2M+03UCEU+rCN5ylzfuUqJSw27KSCkd/
vVPHYv1w1D2F5X9cbyFb8kenHyd5u/+AMwgXskZjcLqWKk3oOAUtYb48mgO8HRRv
W5IAfIwK17jp1Hoe+7ps5B5Mb4XNSrUV6/SDbWxYanUcXhdrZlkwT/T9aOxAJu6O
`protect END_PROTECTED
