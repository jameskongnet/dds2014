`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2QjjkG4hg290zOZh7VAFpo8qD261w5bACXW6k5VVoYK7aoyFnQQOewQ+HXR+Hk84
gkBsh74R1nGiEeW3YmvkzBHflgdxni5QewQRx6xhD411IYpDQkC0L9PRnGScgUJu
A3NQ58PafL+t0agIYzSw8vGQu2MLyr9cKQ73nPQkWI7yWGYfrpk6f+MtIK/p5hDB
mE/2fZbDJTwPrvEB4cKpxPaMYrmDY4xIjuJA3tCb50DDj7jGOr2da7YK0PVrx6SW
Xs6FAS/Sw7eLXcsHDVxu5800oAV1dsqT8jUA7w5NsvTL1WTHlcNKyZcSHWeiPdCa
z6p1WDsWqNYeCBkzJqHbsotNugjHBqecPxlw0N4ZMPYJRnhYEylNQdMVxBrGSrT6
M9mneWDC175Ou57uU1m52DbrLAnYDo5D87bOP2dLCEhEZrzcMJpGNDz664ziUq+0
SjD4aw2s9V8d+i3/CiY89TewBYHrNWlvBXQAX9LU1hUzGJNEmAsT+yUUpm7wITBH
b0e7PbiqTLwsGdf/lP1IzgVTOyEsSrFRt5K5ZKl6Ke2JYxEXFEgltM0xTBv9mxQK
vLmTjAEh3FhdQRRteADo/9+sB+zpRjK2LW969u1vYAkYzVy2Rh2UUDNb6aOtq+RS
ThdKVDQ0ROl9nBKd11sncBFjHlsOnmM8e5uG0dEgZUesJ1EqPAc69+16DgfDPaKL
8hIGgFxBVw06weeX0+leG+oMb4mYqX9kcH5SgFu7aozvzDdMCoO5F6+46bA8yvzx
7F3Y80pszcxNVNfcvipPTT+gu0fCLgpyqzmvAcsJlW2GgCTdFNltrYD4zwJN+W17
`protect END_PROTECTED
