`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4hI4mOZ3UpgFo4/9eaqajrPbhIsmtOhjN0hge6tRnWj8tGm6c2dOom3Cv4LWBmKO
MG/22VkXeRQkZCgiQ34ej63dkUsMGOyPDzPqQuvCh1boTwMyoNTHxsHi7FNafzpZ
lIp9VlMFNAvdLOF0Z3uJQUEiIYbY6h7I/tKwmXteBNjmwXfFcl4JSJVjk+dGNqo9
q4dX467vampmwc+MYjCzvN5mpaIZWgDZQ8sj1kZw4JUUusX2RQ/ixZ54KQ91PZ/K
XyJ9dyiNROpq6101oNBmXgn8ytU9h2V12iDoPAyoNxX/sFqf7T6Cwz6IrnzR2VTn
8TBxz/Tx6gqDJxXxEZqID9nxyagFEcghoiWc+55SvGuBqomKQ5VK2JH7uKalxP1G
HSspa3FGLi80nQUzUpdF7G6c1igyGnpp/XowHS2kxc3ye1MVhV+v0RXDSU+wWJmp
IyRN8/AXA7COATkQ1IQvqVZ2up14xYCuU48+IgMpgIZKvu0C5xFUwRWKQYLpQyZy
CqBkZOuFY0Z+7+2EDd1Rzit4cOMaUO1OcDtPxYYvIQG73l6nsZGdz+RcdHvEsBlW
g/sykROwFovQf4cqha6FVkDxxZn9YkmrBliM2Iapmsg7Kkt7KcxQcHv5OnMXtQDG
e+laAb0QitAOwWSCradzqkYfc68iqh03AUN6BUS2Qrl3pyyWEjNk5F+FK5LM8dq0
Q2VWKWckD0L8FQePvPbfQeoU1z844K4KJiiFSUzV/1EJFTsstdsO15CuzitWhMGS
eVSPvf4bCXTL9qtNEgq7lXLdQhR8azvKR7bgIh3hflsLbbMAoDet+lmV5b9406A+
o16aohDnZvq4vgN5FYtClbKGIEopXKXwEtXvVPwREt6eRByEu8oVuijlSo0/bLmf
0KJoRyrQ7Wuu+thmPPajDTjej9DqiVWqtgbYim4ATftcKysrDk79awWxNLkw89PE
o7qyCzyG7o6gKi7O5SVMJogE2ZZuEd6onxk3vpNUVAK5/0BVtaGCvZV+QQ+siAbW
fG+s+ngHs7mljdIf9eZWlozVT/UlL0fWjAHBMIsxGKwYgZe84ZPW4VrjepmoJUU2
3BbESUgjFvWLFY2QCZ3NX92cNg/WWy4d30l9n+hgA98AbOYfbsOWURAPaf8ogE8c
mXJNjr2Iuf5E4Nrkc+WkZbjSANwYZY08qiPO/ASbifRX4mqHarVuOQP5yFXM1V2Q
XmUF3TMVfOGhr8GLVQvM9WUIhZYUCFFHm+0pPdEFQqS4oAApjR3sjrS3+G+jemSB
qh7I6EcK43mPDVfaLp0iP5a0fR6ogp14CjtAr0k9gZe33amA3758BUXDtMrBQ69X
rDJScdt4cVfZXmak4dftrEXiHE83Gap5LLj5C6qtkstsWFyPqY5uFphxWOksUPnd
BtnSqds+2d8kBtg3o2rrU9Gmdoolb0lKiKB8C98ptvlk0w1CWEynqmZYaXAWWcqQ
KduM6miS1jHH0RRJFYoO3NK0GAvyQjFFmn4lPa0LDGO7lIHeGrjNVM+JJQXr55AC
PvyREkSt1Ixi+1EQKJpgabX3xnMu5omStGtp91dyWzE55KglvfSFaCEfGCSG4eVa
9Vxh9GEUOigiSSI04lmQ7jOhPUHBfE3YOd0avVE5Pzn1vFoDBT15Kw31FfSc1R/q
RD8eOL0z16tgyJUsPdegPWiJPq0L6d6Vb4IwubTyO0PRIkmQEqQpIzNC5lkEoGZ6
YRKg6akxTtyN6bdpIaBJWf66qaIljVshlLnKxjUqCsF6Nd0PQUDNy8jztIqTthXv
GWgFahImrN31EVE6Zbc6En0xSN7GoPsJhuJI+nr1QYNkSKTjTecPi6vngVsGLAuq
sr818wsxcYw6ooN7LHPc++BAwTr7SN18X+D1Jp47xvfstNR2jGwjimqm337+Orvf
3y4fujQz7VZDrl8Qi2Y3hw+0QicY/W4BkZJ7gYYoBoUjJPEbc0YEQDsXtdwPWcLB
Yer51T8gow68JcJ4nBAhkg0ErahmAkoZ6DhTct2IJv9kvsBlhhPyRrJhiR3cdVnx
CgvWQZfU0EtyW21IUgH4Q4Afg7ZjMzh4ECrglS3ACkifE/Zw2GCtwNl+fh+FNQLT
XtbepkpE1wRTa0xKM7igi8jGxp4uo7fVEBudPSXtovFeHO9/DSPf9zFZzf52Zmr+
olJrNZGqYWA9sbIsfM87RdmknfuCL3FBbXxtsk6KT+Mb0adwb1n7yw1SqJJFTOXn
jsYZQtfv0y5KR0+zPALidzR/fuE/GzeyaFN9cuZ17Ts=
`protect END_PROTECTED
