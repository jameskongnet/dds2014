`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cDanyQ36Y+uspMSyliP54zT5C1gElt1uEtcwDI5Q0LYMPeTQrvJuvjceErxwJvbM
SMKow8227IhFKjA8zL+OoyicfNY5ZaYFtMX0Ea274vAif1o7xW7e9UkB+6rx2Pfv
Pv4OsubbGwqvSU4YJYlZZGy/MpwfVrrqmdHm9qtoEJICZzWDuMNcosBR4baCXxph
E0cblEqzWr1NVhZd7Q89x0T3o70LBPZj4XP3Vul3lYK0PG4m1khXWv9HD1yu2iLa
8KVgquwYh03I7tZZyF3LO5g2eT4G86hFrgO/9pUzsD9/FcOA/GCIgL5eE3CFdeJR
nMDdQ9hrSrbTJkM29dIvoa/JsdXEuysXa4OyIJCImDwYVEbBGEQIi57tttOe8o8/
+U/cUnelfohfUN9ZIhLp9VudQ65KvMz/gYroJEu9EWES1e2u63oKh7Xil3xqncoM
8eo2TVpquGVC1IaZzK0GvxO+3ZBxMWByU6Unw95RM+WveTdtnqSHxoZUUdRcCB8B
WqUAijPQoS/dK3euD8Zcab4oDa3WMDse5ufb9YSg/b6ndYIY0bt6YIQVQjgYwuPE
Kf6iqx0EBM1Ir7MbqrN++4NawryNhJiZxrxZQ5aelltwxo7iFGEmDFucP+lln0Tm
/JX3ooRFTAHwE6dQY6D4dDPZicnSku88YqujoAer4lWGu3T9UcLx7DvPVLwz39Rn
cQ6CWGAl7C5rlBosXVaEjf44gmgvkfp2oKnJKmJAl84JuyUPM8i9vqZDslgYQQr/
g18urHYvDo0sEelH1ke/Dxhz2xJc36UiTlV/+o/aNp3tRnceiAT5G/2xyUy+hG8z
vP95GVPHRXkTuh5BOnS9IElZYl81MMV2d1SYa43IZMnDaapw9NCuf/aC8KSzonjV
WqcpA6a7+JUSK8gtcm3SfmRE8+ghuzB92UONwO5OduXa5kEKeMGHhYI0/9s9uYGk
K5K3HGK6LZNDZ6vdMJbGE7aERsajrvKeCKTBRL1UFt8GlEnFB4NNBea+3hSqIT0T
Lf7gCLoTc5JUzfOvUphLzdUc6nS1Kldx5alDLzE5Q9pnCXYimkXsFysBdTCvuXBc
sdEa5OCuWBtGrxMW6fYUasXxtuhL6eIRAWs82uv6Uk6kl4RHrBkpHhAmCW0bROYt
gIZwdIGAP3saqKbNSmyrdhGFHcGGIBhmK/UXm1m0UEj5ifqPxPQpIIc3IhGsVT9D
D8vTX0qtP0/hCnmV8OqLmaYdUxwpGGzJTxIjOm2xjL4=
`protect END_PROTECTED
