`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dnVe9e21W2WHrzNCFhjSAY0nwBlGWn6aLeYEcRxuvDe/a53bpoRC0SSnBt888cAj
CBygg60kMkPPWmiUrlbiNh+oSmkupAlAU7Xb4x0XfZ18Vdx7cLETSA8hicb+96GE
vxy4KIHb/1BNxP1VwNGbAbEHZvjV81qC0fERmUnKEksZzA6pshw6VBaLvF2HsLW+
IinkYYMukQVHFYiv9STlLMtfjp1fA2BdVm8/CInvvSmISjyGF01symmno3h7SQmX
8+whKATkWWWxOC+y74cjnpm0qALI/ma6lW0W/IWqst1iVyjXQi3XRWIcWAm3xZiL
ioICMgruBhUw8Zqv/f0bPjx+AAy5SdOhLekfiG/GExKoBhoD0wWjjyPPWz2VVD1k
2effnyQ9FjmkbqZJLAQUzM+iaaavAiumD5vVtzdvtAQ0A9lfsMVCV6RySGgN+H+P
LvznN8nIo/RB+nsdW/W3da7sKY6ZjamyhqiEQdf97dRckVmdkSBQ77tdF9XZIYen
+Cp/aBMfsuB3lWOdWFv9k+rdFM4dhS+W+7Ij3NLOId5f1itQdoHbWHLORjYj/arT
olniA9qbza24BL69AUtKTJMTopFMowW9YRNUQjAP2gVW/c7x0TW9OCUUodsRZXU+
tiWUF0jU4Lt8gPb4dzXWzu+IDaGTwfMaPq3gYQ7WwU/oihhNJnanmayE/FvZ25HD
R6txlKROOnADc9hybdqCZX0ybd9/VfI+ADf1b7vCgRscBuKpg6KhyPK5jw7S+WIJ
dMah0B5XQ5Rl47b68h1fSQS6RLxRWYblPJYdmb3HhlhWDEBPBao7xX/k70KeaRyx
J3e1RQoRe3yXBNy+zRXmEAQVV2D6KHtrQbfcnT1CsdtZZKEua2O+VwCRDr08wejR
BVP15VrLhJ4y2AH4wquMT5nODrlzl+LGkIF10/Fz9+BmFhIatuFpGErYVcyY7o0T
9htHZMYmos+JIKK91A9xzhg5nymp6Bg14AbaVoRAI4H3CIXmXEEEleqDNIpL0zq3
vMSRDh5mAk8xUqL4ciC8Fxet0DKLLxAteZ3rr3XCLyJfES+m7bagVUk/MV+o3dki
0n3Qskh/K/3xu6yPaoFLIrBTORloSwNM/pSZuNmYEraBVQc4VmMSOGTeyoeoZk6j
fdncwB4yOF1MCD5hCCEX8by+8V0NPgLgCQ1KEXfs/fkrHegI3Y+Ka7MAkSPXEip6
GKYn7truN7jvLOCn8RXqeA==
`protect END_PROTECTED
