// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
WOBV52dk6EBWBs24zMxHl0eC4w8jvPTDZzVsvKFFGnwDIVQVs7wripu9p9VDmaRe2Hep21Wvmc57
8Tc+m9MPYB8i/BTE8wqQIv8WPVWV9GNkjVXH5M+wpU1LBy+DFqGsPbCUDI3CZ/urXMWfpqwU4T6E
9NEnquh+abVrtO7wEoJTAykChpfp0EVbfgGVsnrQvzdB1xsQtDXlCeiOpZg87PcWfdo+aq7rQ55t
deoKU5AOemdwj7anKOnWOHSnUvNAspMeGJkgtWv4Vq6OSHF+lmz3drtQIlNGtIUHrOw2QQtgJum2
dP/bZcNIAlfrFHGGUbOq92jPiYIFVabXA8k5nw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
VNZjhxYhlv5bHPBILDG2ks+PE31ErXoc5aEGws3bfYObdq0FVsN7tWL6WrPTbbif2e2/LopM2eJ4
yMqd3LQFCdGO15Ccn+EjN8YjuelqfaGnOWi4RS1Atq8hY21BeNRLrTdqW1CY5wMD7MvAhVzDIj6D
fEs4zUUR902DGDm45FWuQoVWwlni7G5L1Kf/oHpr3OgmzJdAo8qXV6cKz3tUDNAXz1Ff+/HNr/Ut
XGF3M0hvnCNkFLWA3tzBFr0Szz1aiOcS3ICu9TDDlyfXduvoGtrCezc3yrLQWlJl2e25QUYEiKlO
IRFPt6fobkaDjK2ET0AT6hqOYDyrsuxounFlB75TgQ3z820uyM5wQoRE61aoK9m2y5PeJ3SoBDZb
l6KTqgkgrt4epcdUEjFeYdS0qpMpl98/rCdVDnAe5iRk2HRsemmc9uOpV/rH5EAjsQoENlAl9xcD
h0gOc9Nsr3RJbA6+t2uI31A3CH9CE72iUjJOyU6XjdfbDY6mtQyAMtIyD522Sos02eu1GAQB5Ttf
oNHmFwkV3OnWdL5L6miyLt0MIdr42DG0w8W6l52IC812rRu5DU7sujrishQ7Fmed6Cn8E6zJABD6
qI6zOFWveiyWcWi4DO+dpA1xjKgsEXvCBcCz/Z5uWRhsHbpL2FZh0ripoM8NEvk5owkBXCL6CbfL
I3BwQv9QfX5dCfumrlL65/bq9O/kuvP/gto1wpJE+CT38mI/Ck3imB1/9aa/DNNqTyu9Z8f+xU1t
mNF8IcCqSx6/VwCAV8fRdMNqcrzxXCMUOYf0VOIZe+VuVktlkEb/WBZ3FGutJoTlueC7PeLZQUM3
lpuB4bpnwSY83CiH1vsb2f2tKK5DDcxJwCtDnpfadRk5o7sP0a8917nEuAP0BQyF0/JDPjiUqi2i
HUe9W2YiX/D+uNX9AAWtjrrOf+MGP3iyUtV3y+lgk77syOZyIBd1Gu3MxFOuW8/J7ExvQvNIvKoz
C3ZVpn2ybRMpG0MeTnzxud3MOjfTXBha1argXNeexf++jJRo4LJ0BewbFZ0zIqY1uqpAFx0ZmzVT
H8FB9oX7pXL23NTXINq7o4IaXDKgRRKXDPOB6IS8xLbxqMqJV4x3WE46syMKiYr7ifcOdlIUN7Nw
Gji6/R2OVWH7PW6yZqcoWaMoyiW6H8uYhkS4/vUM0xPzjW20KyUPYkuNWIxiG5RAzlwKNtTCjcrC
mvY/IOSH4jkw0Kjiz3tLD0O83gXo7ZUWBrpKmAEsRTsLWgIxj6ksJASkHC7FWp/YDDW/uFKPl1Xs
tGc1HIT7u91nFwz0XniYxzmFs8TW3zDaH+Qv9WQkeQW7c93bTQTRysT0rnCoPDUxfiUqGZpp/9L7
FaWnPYTkZAs6ZlXMi6FjDFQ20YfC+xFGGNyHI/TZ46uAXBQg2pnzqrr0/eKcc4KY89RLuTI3xVru
xcBZ7KIGbVjuuSR/wPikLYMNQSsGPG11E6M1Qfypy8TvGepvwfbH6kaMVDSUaGzQ5mOHfP4pcmIu
6xzzarE1ei1qWJjIe8sbggQ8KhrLtoITu1vGvcm1S6YH4zk8yWzAdnAVgnsxo1JXVOWMyh9OOM+c
VuElO+DETs2hNS8Tsgl9X+zaxbnwLuvPcwKt1eiQNzOr4GSizyrZzOWj5HHGgKkr9pg7QnBTVMNJ
pxlZ+YuIbbUcgQ2kTQZRmx59fMVnI1+FOEuLBflwDR1jYhwpOx17NLYn+rLNdjqEbX2lrofhxykB
yo55LFez3LR83LITvnIMlEFBKj740Fj1Azyfy2Tn5qCcH8Edn3rboX26e7gaCdetdHzWe0Kqlno4
RvkCMsqoTdwe14yZSh6+Yd9hhaftrMZ8SM3gASk+QSAjaRh3SpP56OI4gI5hrUHCXQEZNHCIB+KW
JO7oS2u0vmacjR6iQ41mAITfqyQLghNYFUNgMRDzEwbltgdlEyirxtheLl37OwHWErkcAQDbNMi7
kApDxwKlaYfj0tOvSjQBAX9+w+wlRIPHBFxP2nSxW9giD+hABT3YgkBOAbKurrU3Fg6QAdXB1nuQ
Ya72cxDqBpcVPb2val/omDyF1FT4YghADI6eQLEYlR2R9yNL5AW1zgsLtNja7stOXLl8OBggv0U8
vKqowGr4m+oFuq/lR0SC2IN9IKumJv2CQFYWObkBb1bJKmHc8icVSy/BZFv3KqpG4SUQi/kfGhHI
xqALJls9ZxKwPqGwxIOsKlf5ak4isXwtnSyxnnABamE+/kvektn9u+7sBRXS/tpR5PXzmCYheDdm
K4xraZ/EFi7kwIKtnGQXUPFuHtaOspUmr5Jczx1G7foRIJTJitVb2vjRm4JZ2oQWHi9xtgDoCJk1
E5d/Pu+OmIm9JtvmrioAjPWGvxJgVSncfdYGZZMYUNyFIzfm+V58dF4O9IZmFAuzJm4xPI+MpEG4
hAiD5Z7jSi+ia1tQisaqBR/83kBKpGowK7ENUTOznuTJb0abiku7MZfJX3+g+TCk4ujCxhIKvqs1
enCQloyu2V1iqRuWZvqYLNwo80dWfQN7x/24HVTauqee8f9SWwr8czMtBFpqo+IWckMpXfjw3dPF
z3V5Bp6MDQcWs2YF+jABALZFkERe+oA20c7CfdkSxCx8dxX59BPmBkSiYjvfDZ9qHtJSoYgewIFf
Fu7wss23zEu7I20WHuz7WKemjgpAjL+nysKvNsJk/0LX2Rm4w9JRLemccYTEMpXDJXpbUNFg6RMe
uYVp59N15ItRFWOoW6SXY4VE6vRUo72JjDK4Tx6p+9woOsrR5LzT9UXaJxIURlPCtFrrb632Tkwe
y/wU9vYd6Xy904/qyDfzhkwHp1b9AtftgEdmOu64Q1I0Yjn37DR5NPtsEZr9YOqiODl/fGmMgSzA
n5j1hZOKSrDf+Ny0Vvu+Q+YKRjYITRaEXlG4NvTdG09ulNh8GAHpfVjYvscSe+WiljRGsLIAT3/O
+Ne4WJ6R9MFz6GF6jr5+NY/yoyoPR/sAbOU9chqgMdTPLo1ezUN5M4aS+FnnhrZhDPAUUQs8aW43
3Px3xS+IMNHEEcVlB4/mtGq/S0qeaGa3b3X61/lp3d8yqn9p0VpE40mVJtb6N9c/699BTeLuB/S1
VOPA/K6OKNf1ETBeOUSXv5PYdxkoZOR79/sgoowkLGvY4a1n8rDkRxDh1Ubu072WO6CZJCFr69Mf
Mahc5e64pmiTzzl5ui5fh8NCO3c/xkSNKGlcFKvu87mYOmLn3SG7AtbIjqRK+1BBHgsFdezCvmnJ
Lv7psYDJO8Ftm5wh1VUVESya5XNtpXuOmxFVmPEcwWBeWSZdO4bu7LJwu56bwP6sm1poRcVTCdjK
lpaydnkgqyOfdX3IfkhAYEgzmxcLdvCsT71WL8L/lfPLKvDaBqaLjnz+apMG9wmf4pB9VpAbAoLo
FsQgTb46LIeORkCfWnQG/MrokyNEV8wnSl4YfFYtyPqatBlA+cgp3keTOCO3wkYMBZDiOTMdrzMx
HoNYA46WdgAdMYinnpg83y9H+NXpXfjd4C8oB6v3Nt2l/QzYTLqXIT0YHRlxSIvmt+rcnVkQo/A3
R8IkFNUEYRW/Ephl3vpfcCNBbReuNp/qx0RCGvN4P1IDNdH6iwcUXv7vqN1d+6Hgxa5hfvIwh+aJ
D8A1NRjkz95aGi4ZFtMXXA5OaG8RM8c3ouTY+sow1mWg/4NZcL9GJgKvdcmAZYuiPgnC6jsOSpAP
qbT1fndtzmZ6ddRdm7/HBRrf2aTmZOHbOfiCMKazifeWcZnfeksUmGVsRZED4X4VPQAkVc+9NHaV
toJ/qiAL1L563lty+Tkt1UTAA830EQa9bPbTxyZ+gnlh71JEnZQdFk2wwdg6gpeugf8nfjNg4rJZ
YsnvZEpInrt0zf9fEbdHdAw3pPYRDTMjGvEozjfze4171htTI4NPKrgma65TdU1ExNB8sHX87XQG
wOnA17WLOzNwIaY/O4QzmvCyeizbqnv93UwhVP/FYfdmgUUKdyVejM9S43HN21ZyIGWGRBtW4NES
fPOvZxh2Wm9bAuNP2PVNe4013UafTWOXYVZ/CysnX9WZGFxWE+BsQw2Q9aace70WQGiQ5TF6BpXM
DtIAPkXBOjSYJSukQLRKi4Wdm2xxxBNMzYuYlKm5vRmvmivUVCW8duElMZqgJADiScrYh63TTi3F
STjhIADnDXJfkYUBC71YLa0p3uzCJcI/0dyczarE3lURO0JlYVxhe/0m3hHx2E5wYTTY+FB9YUWv
K/IpgGSP00ueGWPbKAgsNn2EdXwLcbKyI7RIv2aM1Ur/O1RH/Vxk2jrW4Svg3xEAayVw+hP4UgOI
EwDk12xUYfK3D7plbYoD+3k7KlMlh5wCdmGiaOE9jIqSBKZC9+u0I4cyIO36RZ/zs9h7RhvLP9wG
YS/bRllyk85RU7huxeR/r2Dh+cDq65jd0EJ/qQrE38KgWP+6qgLpS6R5+ygyb+RDqFUQSu/JxIUH
SPQSyYPG6j7zK9c0u22DeQq6BdTEW4+zB1atTVDsK404TD8l1LL786smI+7MDPa74XU7XFIfieWP
sL3ugxQRRwl/JTvfgx//qHmndxveT3EyoWtw6e1tbWaaHzn7UAoUFcLdXpVGBzIFT8yfvBqjaE4r
aV+nZ1+NQxUo/qnqrJY66MUy1lqEItg8m5wF9pqpp06kNMukaSA+fKTa1BBjqIqNvi+bQVkuPAlE
qf34Tdj/be/NO//iu7KHKlAKaLl2eLyRci56jvh0M1QZUnog6Z6WTMh5ui0lZsrs2ILlDHlLrcr0
4sE5lZfe3BgpJZn99Bfr6T0B36JxtnG32SBDRiV9KL/KkXyS4G0JoOgesQ5PXfY8jUfBe141egPS
Y+l+ecAiGQO4tToVL0Zrj0E0sfklZsyTSg8P6Ml5iKD71MIPsMdWL74fH1SwslCDp+MxsTgAHiUD
tMGd937wKlKvtav1uhp8dCRyZCICzYnwNPUAj2HNKmLoAc01rRUNG6I93huFHabJ3B+8eoIme0CH
da06R4ibvtmpZ8CnD8ixkrSDKGyw/ZY1ugJZS0GMnhQ0vbdRn+txZmXGior7O6aVaE8ZDPOKCLdt
pSNvXRRQedzjHMNTRfjRque0ucV0e1E6jVJa4EFyF1NYDuweC/Pv1UaHwreFbTbIKouUD/mb8RrD
lopyjTwoJ8Q/dbp4ve8HkR0bJbs5RlAz1nj7/qlUYzA4WyV6tddFyrw9Of0e2olmV6Q8nS360weR
Drj0ipBYObkVxrUscOVSomeZrGYLfC1d8y5vAMmrBqZWGfcxCp97Zm6zG3oIKXa1Au7rNGVWO+wf
lozlVsG1hMwDU5GoWXjtMmjTqK3IMunl1TBYo0SgUlIZKqQyFxwyLXbJyBxLvKpF9CwwRm3cwn97
PVi+ixGbwgs2wfcJenkZA3sU1aGroAF1vLP2tB3UTJKZms2yuCtJ1yl6usOBOv+7YkKriiSpYGaV
L9SqfG5dmwykA2bTDfhrte3S8jIqf6AjUUWdXDvBi5LFvZPSIIIrmk1rL1yB+OGMNmIjv3aUTZh2
FulSo2QvEejOZpV68TEG5dWo7b6hNQGGkMb/BArHe0dQtit6DyXCfG/17wjelBbdYML3T2cw/TzG
Tpz1IGS1AZ/ar8Nm8Jk4IlJx6eTEzz7vGcLQat3Th/W3rbXB0rp8nmbYdUlhUwkUZVsZYSmqAsnM
RIx9DQVxGCgiGUlpKRRyoqFTzmmyJQWKS/8yfXSiHIApYK/4id6sYv0NDrTmUXg9o+VFkLGHhmBj
6T7MsXOfmBZ7PirNPrXhlNtEnWTWPXoqbULJmRc4ZfVOtNJIJq1+LUB5xx8JuxLDZZWd1tzcjWNc
uL0ldLhTnSgN/bWrnK5uBH3sQyJ0A0PpANIsWsdlbyUnAeCkB+WbnDo6poaKitAksf5h12KFGGuq
Ge5W41M6ckbsdTkHZ1aMUyNoKIX962C2XzCzwVlyBDtu4rIb80hjX0hWTZa9oRB7vpKjiYH9ge3+
o1i3cg12qU9Mm2RDiphXn5IgMTx1BGAEFFFD7wFkd/cQU6OcBTF9QE7DykiCPjhC73oeR6fJRd24
t+tiltwn1ohhaQC76r+sIfjZ84eEWEMgM/EiFQWaAzJhbtWrdCLIjAz8eG7g4fIWP4rxfPY34Ksq
MqvPotimYBzKotRFRh4hF8LS6sL5Sr70foaayBEGWwDS13UhFkMkdgtRXCCaA9H/qlgV5ioUv4k1
OPAvgawwRlK64quBpsKb3RTVkJ1NlDE/UlFHk1RZR/rseRNL7CM1jZJUJNlCtNdtJMF5KJPU2XkG
ViqUaHlqW47R/B05v7NE6/hKaM4ZATtFL90cvQapMfvMGLqyFUK+re/XlcKt7JSuEdjkoB1yWx9G
oTr/clEMzwn7gTWxKAB0NhpikrOCYDe7PQr6tYZLXYsHnu1s/v8uwcDGk8l3HAZ8i9k0S4GPn20v
oYApJmuefp7PE7qK9esy07e28y9e1a4Pd1laFYBhChEpbytdAyMVvJot8CnJi4KBB9Ov/Q12lwcN
g+n8au/tVIDkhme10O9Zn9P/03NA2Ug5L8qLzIDWiuCJji604eGgs7ls1HVbY0M9RTyCoE8Voa+u
c3fJJB6BgS5lBZ4oBniA3bdqh55402hfSsSsop8su5PhNFa5QuceTXaonZveYvE3qZA1ojTMQmW8
E/jmEv9DSNpsq8ErC3hIBCmU09IkF6XL0Cswm+2/OFgD8h+wvgOs/xkuABuffz88ngG32cLkOyxN
K0BUKGn9OA1AgXe1fxbMQgbnzTNw8ha+MxvXsnln/1Own4682+3nmb3TIvqE/lEi9R/6uFKGPao2
G/5kx93/5JOBEYoo6yYlqT7GubwhUfKt58XWTbnn1MOeJ2XD/YmtqPP1wnKaNKwCTpcOXJypu+tE
TrNZmTjLrAcfXtjrL/moBXTD8F5Zlh4DaYvQDixoj/wu298X7IzYVphCDgtqDO70FVjePhShLisJ
sWfCmlbA8dRYvTsla5a/fSztSSwlDIlc3aOrCYXV32FkXV13BcuEU92SMRO5AMQqdApNK/Z5hlHN
Jm8qv1OrOFilir2tORLK76RNq4dSiS0fOEA1IvcTXy71sY6AlIuhiwUXZywmCbCy7Lzun86l3WYA
o7N0nHvVldUrFW3RbXjtJ4Janyd542QDmD5/Oq9QJkh9bNtF8LTGEiTUFZpb7tmaCMlvzTM22qFl
NX8RQp5DKDezbuuq3vUMAz7qC8k7jjoMdvG852gwB/bAn2hhvgNG1/3GielUC/pnp+843xtCiYCI
qW908ds1fAlRzuF41nVhgZub5aOx+bCcluICINtq2qGlFHmBbu772MsFOI1cXphzT1XQVcU+qOnJ
Bau6PpZT0jenREzbzAvlSGs37O/jvjWGm8/l8QypPR24Sir1XUxIJEcquvLr89lZy9wZZjRUMW/r
F+Eq+lE6tk8pzbNeNC6G9kzkIEYuK/xv4COIia4tXHjMlyA+tsWv9ZdAk1pWGqD6qaqwdUCB4UFI
j57fAv/0/bTASg7aVOiGPF5rsXnGgiseUhz95bsBIzYUlSGNlMr80gm30RDI8Yp3OC8u58IsQK84
4SecGBOloujUAXBjLvPjL1C8l4we893whi9Y0Gc6JwV1nVwofmnGYogdN15QWiTZSaAQe9+6bM1n
ysOmZjusXTITzmr5zF+mG8Oyzf4kYa9A/diV8ztP8zAIAZJrszREDb6lJi5WOh7JuBmupa5t1zNC
VUq3+2kLvYIn1TtQsrXoAtIDm+Xs1reliWuuoit3PQeg1kDQcfa7AS08zzcMLY+NQ0A6h3hSHmHu
5AlL8VUx3c6T8BydrA2eWptAmmjhwOWq88QJTBG2cAREHtwLo5gndBS237dgpfpa2lPXw6KDmGdL
hiobATolVKDP5egoody8sv14zMDvlCvVQ8A2S0o0o5u6fxt6XVJDXufavfz7zqLiQoR6vSrkuZYe
tsDm4r6qkr3UlnkdWj3MCAiR/ORHLcrL1+8rvRskKJIAzMee/48r4gtT+/g0ZYoUSTKKGLMq8jHq
sDyVaLoQ1ewfEzWYPKVxc04Lpu8pk6fvRmPie5yMUXq475GlppBiwzSxXuJAzeFjZixW3CA+vZuH
We7UDjaWD7v4u5JJ1+HQZ7LpkKD7S+2t2l+/CozbS4xPQFGyfQUhaCMtgdm6u1HIi0LajzN8fBRj
OYgemgkG+qgXXeH+ti9Pzl7OC0QIfCmSpY608RvHn+66qzbqd1sZC8As0zosVroWA7r6gtoRQaf+
3YnKQCgc2tnrMHiLRBVTlFoUBKIJ3/44avLAZP/xaEgt/DV9XMCAaOLZrDeeptOeH9QIDyu3tsiI
MmJxVJYG7XSTtPIcM9tMS78WqtjOo0xpVZMyYnb5dwjVWbAz6qa70dJOv3dtjeovPEqpn/oHuqU2
YyfvTchBjM5f
`pragma protect end_protected
