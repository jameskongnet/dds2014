`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9BmRbafCgDeUopFFc4398gXk51gzbfr21GQmOy0Zchjpp61to9e6QlCCK6+rEkLT
0kDBioMbYeIt7Qq27/j88//ySOQNuPueq3rabNjC2fk9o/TDdZTPpbAXiGgDosQD
V/UM4IgSo/Er5kvYS6KOHMorSxwAxX3n6ToZrZkJ1AxK9qb6CJfxVVgM/kMx3+60
E60V5XvYHfUoSHVOtFhtL87BLrHncFESKbspYLw6LQ7FVRSF/69H0/9Wl4TTjYT7
VSG4fIy9hOGq+6tQzntFa1rLcQJe9O+buHUCTVNS2Uzz6buahQpVEzBA8BepODqM
IO4xsQ7b4zBn3d/dR6Ocsp3rx7GPoP49AgGmmXBpzV4DFqvhP7w+/GHGhs78NRa9
iZEceFsZRR3h7dVl/dBJ9bhwvsApQ6gaPG5F+38gRIcxXdNGwQgUvVLhCuXJI/2r
KT6H5IMxuCcky/G9+jvUu9QYkI60o4uPJr7FnQ/tHSBUK31/PTwPSlsh4tuWFk9V
cHPzvMX5g0WkknFhH544mueGaCDNh3h3DDUQJVLo0nylO5gdlFjwHstJxKKZ+m1s
eop5iQsu/RXCDUc4i6lIPZBBMaY+lbHzxiCqD41bAO9IfZRaMXzeZogLhpa787Ry
9P8h3hmUyJYiO3d/Sbdtxy2yTXPGHUDfF07hy83VrDYt9ttvpcqrgWScSOOmc4G2
ZMYh1+4BvQYwq/StZNSHkpf39RP3QpAxD0pscaZS+FWRFPaSsUkkzI3mgFGkevFn
tqhG6+gJKC12khVsXG4zOMRc3T2AjOF/zWixzub7wEZuLvIMveXiT3R1dmLMFUPq
tbQZceIANrmDH8J8j93j5Z+UjIvUXdEbnnHkLPeEk9vMmvD6p+buy4roveJFu+zY
Ajek+hszQ3T+lBjiBRXh+ZsTrx+jtBl9FeR5ZJDoT1+OD6FH98v5G0JiMaoKaGeO
wByXeerthX7vLbpORhdztwyap6WFFJlW+70zkffqNKcu9Nq8rLP6lxPZbzwTdBIC
3U5wVoo6x/DwS+rSYUM6iBS7tEFJwFTm9kBcDeswWiQavaI7HgaAYn1vwFHzlLZb
InA6mGYiU8mQxLQo+58+jsAz9hE3uG4fXlYLfj/lI0s2OxUnaUicIIx+IT3ga1L3
uM0mWhMEYZo3XGiEmHnSjGX3DdqegKg1/zPTPwi/wt6f1SxmGenxThjia6phXyIv
JDihv863ztuwmE5ad1aUJO+CYN2UgVGe27kd6onjpo1p5Zqu8x8bujRffpIL3BuW
97vkaa7l2iimh+ExZBlU55CKtK7dh+FmSqMzvLs6nOAAHvXm9BNjZkXIhYhqjdMe
CM1qULRTWVNGKb+5uL+ZXv3UWNaikDEsHwkZCwqf4WU=
`protect END_PROTECTED
