`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZKPvVcYy+nXnO35O3i1oTDRIl2xSHeTuupyFS+8CfYAIbfdqvRCdt4Gq1t9OMSaA
mxCy+3Tn9thP4pRyHCCJyFQyDD+5SKpGroTebqfPX2ka6iY8ViY5Rw4/B83HPKOA
W+Hr9nTi0Xju6Dx8b77SZqfnl4BORa2J7NmvFF8Cpjg/lDc/UDkDMMpDyJ+8YIAW
bg183nUk7D4Lmvl0j9GwAg9P7hJtEvc5rRl+lHYOqZYb1eBOvekz4/55E9R39w/w
j+SZB/WdbO6/0esKuZtnYJMe1Lp2I58MbrNg5bFNFj7hk3VQ2tVYIbwfX7EEqrWH
Jr788y0nLABbVySTCNQ26BLSbWI4hnbSR/afbhma8WVERcbEpF4CovWQJNSILRQu
1GfXBi/rQXK6rXOrrdWuuoM1Kam72g2Dwou48dAjAc34TJ1tDh+PawsbLyKCw4mr
esQ6R0DWPBoI6bSrboFr7dMTIduQQAu5IdwxR4u37kPbxq5G4dCsVxihdFYrfdJU
xFBSGvR2paZQIz4d5OwFTUNVSMCo2In8mdIBG1YoNr2zAZfnJA+jpZM23MRds+nh
ecBaR7WZCnYRrIuQMa8qBXwr86+1i3Z0bwJf8v4NxGIgifyi3PQj0RVpwYM4zHBs
Q4C+aMEgkVGOqYO+vVvge/AhTMjVhe4cXOzoKzOoi21AFgYjIX9pX5xDkjyyr3xr
jW9wVWvBtsJIzUuiDaqlrriNJyFnNrrbLW2QU/Y8mNKH3RiILY7HaoEcKDD8DtZn
PLMgdZ0O2CopQtRk12QLxL4bp4xPUpU2/pLuyRBsS672mkJSdP2f+PDkg/0TOlz2
L3HxSA3n3MXVNUfuMLzSSMnAE6LeuxapVPPyIR3evFGoxPrkLjtTm3JcYEQAAS0E
xRs0B9BmzggXonyl792PEeLNxFMzAIa5jLENyf4geHabrrktIAgyVYbj543xedaV
r68EZKVS77YPuhv9H+62nqxsXB3FovsL3wzg4Wsf7I4nHFDx2dmQrBEYgUripSfX
I0vwlzXfEbBKWaTz1TU2C2YRYps8lYtnc8POsQqKcnukd8fgh3ftKa4dKOi1CCcK
F9Zv6Ptjz5ppm1PNXqddIK0LQOoT4G93oajpTl3A15B6M1Av/+eke98p0jdoMGLM
pptHUvcHQYuSz8hSJ+JeBjmApbTxu5taqCqqJ5S+jLOturP9B37yVp17h5+qUseq
VIVaMWTYa6au1B7l15nQkalEmkavMHIOS0ErI56eWdcJXdOnxUm/bElz5y1SWJeg
JLZyOwijwuj5+BNVxiiCY56sCH5PfrqEWSNy8pUu9Ot+XfCNqyUSuUsek1eOE+oQ
cJozVBi41S9ty3qaPB4IJMHGZh6qUPW1PHD8nQVoS0AJ/0u+GxPNXtZoLRsR1PM2
VqmcOpWKcimfnqq6bS3pltkxg0bkgwEcEE//W7ux4GIEg74wzGExIRZD+LTfONDB
Tv4kBVUeLUVpRx51vUGlZ6K9VjA0XNDxCf3iJlKQw0DyF82gV4SLy8CjMOX65nSV
Bd/o8FTpK31akkM/FVWtQCvuRkenpk5zQ0fwtSwP/axNqeBOrR0Qkq8zd2bldwAm
4CzbGYjBSWsf38+LFDblpGwOoDoBcmQzSPaLKUgnpX4/yH6aCDDsZS334k004fP3
hsGSRDvywaRRa8gH81y9E4Tiuh46Pg6A0J+/iDZHGS/lgE18THv+noC5DQezUnrt
Rc2Y5rM9H8UYBeped0xyMZsG5nJn7Tu5h07AmSXmFknYDr/STTJmivsO5zvlr+WW
UkhJQbaFcRaiSpXsSUh3ppwnWgO61p5EbDCRM4vHC4QwyY9wLUQnGeKl8vcJku6r
CJQZkynzy7qst0x3mcM6GFqS3Ct4Sy5Caf7p9Ww4UjL3AXMYRNGxmy7Qwmpm7GoY
24rD/1ToKXS4PvjqgRuLXr9BZ0mX60Ms7JyAoYvMSMkqdcZYdw/hTXkklmthRIxd
+kLKaf5KCkO+U+BJp3g9vNvQgXVNiZGA3EVX6AwFkqYpNQp4tCOgvmdIb4No1/4j
UsunGMrvNSOE7yO+yJ4H6Xp2oWeQn89mxrkhKgnWEYLIRlaslaQrL4FRssgrHTVY
Oa4ht0/g0Xt8ix5Hj77H6pzMJ+V5lfaNR5dwEXeAAQ2AsKfz+d+ryd4uFgnMVCOC
TnGmhnnEJoNqg7S6th4Z1jpzAWrqgJT0jae1of3qpq5d0opY7NmigX8ntB6c1VM8
GGYK8xmOYOy0YNukksncVOGoWEBUQ9oayePiEbOK70GrjrPqL4gkkCqySrbws5kC
wTOjFkOSTQVfEJ8mpNvx6kOXTOQwpBDhWE0DpfXJMMTPTcGTL0rdifrUFX0FwaAz
HAOVpfyi/+/D3rfMyIfsgE7Gj7KlOXJ6709r3DdWhWIx7SmepY/c+/AORA2CPuDJ
50gXoeRgkssz14+TJRiVfslX8TMmhYf8W2UEZwi/Sut3+/RMd5mnblCjmGrEwARG
CnNAPIf+/7/7xD5fP9O94gSixDISYcz+s8SfMfd0d1We50kcRf7TaHXVb7tjyM1y
Vg07fnhWZLuLROCoYxilLkN2fXxUdyx+irIabKntnzloPNBENCBDC8EYKo6ZIVSB
5vGpKyZQM4aHuQPU5hNWGgZbVj2kncmx8zxYu8lZGEQ=
`protect END_PROTECTED
