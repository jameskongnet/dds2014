`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrOqJDDpIbRYJaNMqU4Avhbd4ckbDI5m+MpAvMmHRr2qqILAMmYNcEl7tNt30+Uk
9O0AWSm2CJx2ejkxcU6Hyj9vsTYNZwjhBr0flmVogGY2I4NxLr8g0onMxW3Z0mIF
y5ymjltqYko2hQ8mAcCFj/qOkTo3HGnADvps+BYUOylTPpykdmWZqsRU0rKPyTc9
9+wAjLIx9xdgP7b33ndDmwp7cVsR7vBr4UyqChA6fkR2DONGeiTAUoqSqDLLHCd5
9xVK/5rIgpws7MKPPpdgtoFBlieo1naTnPf14eJKus9DrI98pHm1+ZvFy3N5mYY1
ohemxxW1EhfI4gCUd/NU4cSwiJ4tK+ph4uHL9btECQzCvcm79q7dGcmyZGbZ6H/b
aEaDZUfxIGyJCj+LDzRol0xvNrD8GF+iwN5qnHzIeep4ULUB99II6BGUQAnA2Ie7
7gGMTOuiqv2pF+QlPJK4X+KulgXyd7STMycP8Bh6MWbPyWud7GW/dhjzsAK8zbS+
OH3+x8UoPkN/RAULuTIHL4k61p4l+1MkwKNwnJI4j0Nxmv9Jyws1szJ7Ud3ZwklE
hTPg7NTt27sZvf1TYw+VKQLMrOTtFZZh6qlYOODFSGxXF1ZBR1bFtF/OZFcrc+Oc
blBV75xpmwg3rutBcDBkFFBnT5bnblV6IWnEL39ypJvK8+U3bwbQnF+45eablMkL
tisuHSzKkJml2osNT+/J1PbDXYfanBvKCiHpYMwT+OMvvr1LGumoq/sOItv+cpMW
UMx53NsG2dbWRL6vMBmRtrJ73elEBmDM50zBNXioSB9gAiDti2vcA60bmmUHzWLP
wa+4EdURKeYCiMicXY8cnFUA35QnAAy0gop9b60j7s/T7/3A07ptfB+lzlfiw9QS
h8Gysb2hFtiFF9VbZGe2pKh3xkc3fOq+Dpv+95I7juorTiEvdYbY1hUdWN9zMfG5
wrN6JyvOiqKogZxzw2XcdYUT+ZAZMNfDaL21nHzNfga1/vZop2Q/74mXEmRffKRH
euyDD8miu6XqCX8pRUkhjPvRzP7XoxOM07EYAuRxI/pM9jniLiv3JEzHyfqgG39C
/zGq1dqOSOr0IgJ8WRu13VOb7DQVEMBZS2SrTctDukkkL3EOYhu9ytj4vVf0uo2A
LEDYU4QfXkyLGAOmkeKKwK7TH5FeibE7Yy6e4WOrULB+raoh+aYHW6T2JjoThuSH
0TPf2S7zmByS9Ky99n6xDirQETXU5U8RUxdzRi2zfGwiPnP83doFxLUzhTEuxnIo
D60ABPL2MeoW2uMjAnjgStmYzyHL/ePmSv5WThaHZxn6uLpcyCr9bNIBYuRbQDwy
WVEOdI4RnbDw14kZzoDADeH2OtcCXzZVSX7+aK5y7LRMNUprD60wdkNZzhlOvbaZ
BFsh/VQNPAjEcLGqO5Mt6pi8SArX+Nev3Ldntr4VCKmAALckiTJPkfNHBfg1KCZv
b+1YWQAScm69Q4AAg3ss6mgxJYrbTnOmXetyOyGeo/YyU8H6URHAGSWBFSCrzNt1
GrMetW3BhZxFVSA5rNA+9sgW1ToIU3DUH91JSg8+s9D5VvdBMnlclqrsEdJAxvL9
cC/jfHKbUcBkaKIxJ5sEhdoOu2mF4OHmZkX6sW/hyJEvxOE0hk3UCg36zsiTkf+t
r9GvdIy5Acuc5qFDN4TW//s4w7Zclbb3X/dtKqSqP8kUQE0wfvpzCuk+bIZ5GuOE
UCaEUTKh0weofV57y6MHI2FC5vfp/3uUrzSy5XIxVsU87wW1kaMS/9qqDE0D97am
ZU1jkhQ7c/bpgGlgKQ1waHCS6Vnmq1/bnLMY0v1aP1PByvMIuNGMEKiQDB6XwsTk
fcn+XhXlWrj9zwdm6hWEsu9iiUwVGYybScdr300N9/tKtqKjyV1PrvanE2VqO1SY
iIgoFpO4PBE0ZTgBeyiWHIX1t8cUbNR1ufptGUnQ50eraV3YTDZYp0cszFqGssIE
fOhGGjPDg99PGmNwGINrykxZ7/6RybvVsOokM7Qu3QsKwRhSh8aT2NDKa2FQwICO
QT8waIrNU30sMIRbv3ZJGCt2XXBHGk9aQCpmM5wB3K596aaSVywnrG4t8Vz7B3S1
SoJGryonDO01aJnyYT3Xk30NVwUZizqg2gZS3nQzliVqYQeAEgWyDD1D+vfixOWb
r0fQlmR91yWAUdiuB/rDMlvN2gno1/xKZWwza2zdbLuS4T8bIzYGKqk7fnAzBtKX
clT3shbGtRfo4K88Gp/JZUhCKUCoFtBpUt07l5mc+I7mZ5m7tX3jsskMk0aMmO8L
SOWSO0uLvFumqTbFOU9Wi8a+WX2e9maBDsUz70tJi9Ck2f/+DTrNeRDA+4esNY6R
S8zJeE3FHtOhTrTIYzE9L0nsX9UvT7N04jAGJZeYAujVLMZWg57gRX8Pp5ewuy2g
/TeKwwzyQ4yLy3GfZENbl+cYrK/gfWgL2xsOYDj4HEZqCQn9JCXf8wlKGJhwI/1A
Q5MZ8KjBxmsg+LyKrefmNcRel2eVBbtyzILdIr8FxFd/8twPUNNBEJivh/iOwDmy
HwQg5bUlqOjYl4+wbAxEFD7vrPsNdeP/7oqZ1qSvUbH7/xRcHRSpqEzmbKJTWQOP
IO/D+IRjMT16dATuQsfv83+vXHTCEPoX8qYHlBDli8JPZ2O2Q+1BwbcGRtYJwIzW
9SDAANssmEsyM6jIDUtp+Kctu57U7pMMfGs1yKrFvfI20PeLeerPxR9GV1myvC4L
XiBIrvvMEcWmKyKgOWo3g0sLcTjQtqORup+JVjJwFtz4uiblu1/stFYhvotnqjsn
Hqc62KPXrCRU/3th6zqHCE21l7iInfouW8zTNk3RCqCsnuiVvvjjjdHsbPpNavmm
Msb5pclTrZErejDsDtx0W00xnRvTuZsBuHLnvJ215tefBH9lLQTQrvVcY3s1aNQg
qFIr6XW5Ujvubrlwq1z8mZfdqPE31BaKIuxayxB7nhXpQVsbxs1YDjBJahTEdlfT
y3vLRIwDDahA8mwRJMA/wbEsc2NyXDvGy7/l+7OXDHABYl/zWfN3w/mLmEzZu1LE
ibprO9+x26StgReO+z2bxlnjkFhHfpiroXn891K9BXFxEleGtAjzN8TaLO8oEFxI
Khbqi4ogseQMlyXUvZbW/kTP1yjKnb6E9VbWd+cBIwBUmZTAtRXGdwz+tQQAyC2I
uSKyX969aYiYcY08gMSS4R5u1ccEhQ6jUXPXdHGTQimugUKqHQXCtNB5wAeu0eY1
c8wQXLE8aQqS7DYp+0v7lwvwLVVpbsibDb8p9bk6NJqZk6aY3gqBhbsi+ZlLfkUJ
oIoCTB9+LVgcH6x9t7ptxPA5Ry9Y1rt2Z7BbPYol6Or/yPs7lYEI3NknPFI9M+Wj
0Ep7rRGHVkeUJPiQ5Az9OeanvPYCLZkstUE5Z0TAgI1xFebxrXTZlH5/f1LY0C4Q
TQBjR3giGkLBOYeJfzxOlzrzH9rNbPmAKkkuBRCLzkvyiHl1UGSt4OL+Nh+L7+ex
1MS5440r1hcnRaBldiFB0rYsrgQFnO5cOGDqOL35Qpfg8GELTlWEce6YlAo8HEDo
hXLjQ7FPs/Oiaw8a+OWztjuii454cpQj2VRnU4slP4fCNWsEp8hsSv/oWYcCz7rX
SSGnCKrgQcS5dYbAJgFHrpRJcGGQD/ILeVb2yUttf8n5qJEVVd/buBg7AmKZo3ZV
23Dzy963hAPaESkgVSPThHcpiy3BJB8DiCS8X3tDJ0Zs5vZqXvYDuD+pv/KGP2bU
nkt9oeOn4iDKyUwZanoP9GuXmuUGLbD3jIB1XX8/KwXf/sWzIkb9yd6E//IB18We
/5jyzcYWgPJW8AbmwcEr8kZqmYNfkODrwar+JBOtD+byyODs8EQnBVnHh8QaJSNu
u7yAnlIXH6SobVZ8VTujBn2u++i4hSh8ApGgJYL5wraWKO6x+8nM9vV+w8HLNoPp
zbomKjRwqUgBIP7bsPMZbgCnPUtWcCzbwFRJtPCqt23U1TUbu0ZRk5kZfS6FV0W/
iSCaUChEVn8oNY9kWnryu8GAwNBKO++wKDHRmfxr5NCaMcCtCZ81InnlMwvfB9Zv
WUnBBwNs6xCRwPkWyijBJp8wn0gbxnWJEe+M8932skdGZK/dFgqj9PylcmJLlKxj
0ZDdlypxnZbmVekFL6dPQmAWmGhKo9Sw3KXBfG0+9vQnVcp6JuFTRTcLS50ewCme
lJrcVJBvA0SA3Bk4ZIc9cQoYqM4O5YAe/7DUy8FCzpJJjhY24B/GoLmQycBgXDEi
tTVhDSGrKmNeooHVHC9m99PiCyGJ01qriY9Bl0mPwgBXVGSu4szLVSJLu1ZjePps
OaPgdntmQFJL/e0o7NzRQmurkYpB5xPMg5+5EJ/rVYCn/qy3Ljvz3zcQQFk7derw
axJSEpwj+h7QeFn9h/IzWjHgUW73EFgLyAiYc0DElL7m24/Od05Rg1XFTGPcKyJz
4/NjgDii7BnbrH8YzME6lr4+KoP7KMbsgQ4jKQksnYaNfXiuqEKymdOBLZlLcLlB
DMFLXbFBK3Bq6gl3PeTTqEOaU44ekfX2yx4luAr4ge5uKUxnwrOGhjZUaTwg1+hn
En5WMfGihFjGkfpy38RimyJPCF5emXDfz9dOBiqXjaQcRXQnjFMqUGMMKPKawxiY
sbwa3iVlUKo25gddXC7t8tdVsaNbR+B5w05hcSzTQKeNN3fr+wuhswxptgWZIgHc
B8XTLF8/wWfasjIsLaN7KJs1W5PCmCrUGWgK/ytybAIv7/jfs8msoZjpKHWTkkrR
72txxhy6cVckT3HhQ7o1rJeNrC8vc0IPJ8FA2LhHUNzMj4dqUZp2SH8U+DiO7T1K
SDUY/7285Gr+kcYVWs1F6ZdXBWgyMjc0vPeqQ2wa4sdwt49h4l7twJ9iv7cvQaRG
XQGoF68+KfAkkAVAQhCE77/VmEsN7bYvlc17LfSSyxx/CBPjCpwfFghWUQk/epFw
3Nu8glo8qoaJhsTe9PAng0mJ7bGa6lgEZaKllfqPjlW7T9/bk1E1KiXNyLekdR3e
lFQMe6S/DqDDzxkQOD+A3fICfdZn6X1SiY34gjRsqzjJwE98Y5BxlnG7S7w6CtGO
OI84G2TVYdkpcnoWAc6ynAz4Qx/cMA33MuyCARBSdU2W38muTwDe0uXLL+3ZbGja
LzKHr/qV9KTPgjjD7b2dzk9hbTZoqJfwAj+cw4JB5nTeJWrNw2ha4+08Y3e33Mul
pa4CEN4E9623WjAPQiY9MAD0r+RscJHtejZhzlpxeAQ7I2mpQe4WzN7xQoeYZ0fp
Orv4ZzTI34/vi4+yK7+20fV2ph5dlC1g4+4/5wdBqT3TLtCJPt6ysRbKk5g5e+vF
86V1AnH+dj9Kq7pwEa9cEi4CJoSevWNkGIjqqnlTCaxXS+zFaQEe7a+MDmZBURyg
1pX2V9feRsK+Oidz/FCI/mA8nJ13c77Yk/KRhHMlIfq8yypr5M0trOZa5uDiBHBY
/4yYPDLdC41G6jgEtahknAe5zTIOGKPEspjgSuqJMDMCQJ0I1TNIt/33DehXBV6O
gRkPocR6VQPv72vfWY2UBuaXxVje4Whik5Vfg3SEA+wd3k2GgLiuw9G+XCV1WYmE
UkqsMronGugcj+QK3SxxAfS5v0+VVKqCKjdCl0M0NpK8yqU2U5vanuELckI1Dvgg
FDc+YHgHZqOve2nbToM0Dwl+qqWeTTW42IVrYGZ3qU0FM5rTrPFzsfnkJsi8O6JK
8pxsr03RZwRgKaaag5JlXF63jY58jJ85oyTCU5Enk1seJ7q8+JnlTIJADq+ndvaa
w3xUEfzZ0e+4LFsaRQvnAEx6WwGPjDcFs3JWWDl8t/C7Yy6GHXJE1RpfxQY/pAfv
NBlr1Hd0ROI0dBPK95OEls8RRG7Tp17zFP2e9iKyXkzg4rjmTJtAQKD2+kUjRdEJ
4v622sV5V848gK/25r26lx3AIyWuWBWxyXrHZ7YTatIfq43TqMMHmYCVneWcHWuG
313kOzYVbUe7FrftZXz5IZnAU6HcNslYS7+DhD0F1N++j8uYlBCitcqLW1cyaNkV
YoVuyoqqXQ/MwVCzVrXAxUFm5xZaR4PDG+i/ZnMIZvUeg2cwypRG6OM+jiP0rPhx
5gzP1EE53tWvc9/XZQxd2yPyq7Ia1Xfa1CvSCoHVY6o7avj5ovC/3LzeosA7uh4w
eJ1Pqq1CSULKsk4hdmgK+jzC4Y4Bmb76kCo3c5hheRZSDR4QDXDnvGCygFg0WIKE
YA9Ff8ROD2F0yloes4GCr2+wvprcOG9NwJSF47jtkdx+UUNdUQZ5qMTqBa2LKSFN
/wGWDNqfnyXkikOO80dY+8Jd85Y2Zw8yrBQk/gknO3F9h3gvqkIvF1hzugUYT79h
ZGdmJYgVVIHKbp5cv+NUkQB0o9p6tDwVYkureLvXze7/eItLsykW1yI4ZGhUNn+m
QNEPzchtNnq2gBBOyN8fn4+gNnp1TahkchIK9P8/cZ/6RZi5aEBchvIqyMgG17A9
mTu7kmHE1PXAWR0d2fuarqSXSjyaJT85UbhSfZkCszL8WlKNtldWgGes8CJ+WkHv
2eNwV9ICTMqKBmUKLhXy6XqQTTdETma74PsHaHyvAKvUOwfXE9s4FR0pe8xEF2ii
O0CKzUGpUWJztfQc0OK8xFYV2lEhsrFFnvcUYDav/jnvDpKL6PHZPGS6zfiBAkVi
mO7h4/KW2SsX0YcIDhkD6pS5h0+4zOYx9jVGs+MKBPMdR7rHSSOdPrxmsq7cIF89
eIOLW7+PVBRH/2mlXuMVeGKUlV9KUxFDE/riYdZkbtLsWHNCMdV07VpgqZ8WWrHw
WpnK/S60yoMCSgCfj1+8wMEFCjnom2q/uCChDc7TsaOWcVu1LqVFFCJf83hQazkr
NlHVHLL4Wv0TKbhg2KeRxD/G9eDM48fboQeEviuwUvhPJJoZgqazklO3FvjB1NX2
zjkSZPVNf9e3mbRPI3XccbmG48uCYvmM9NhOgZdvbJx4ZHlyxci0IUscAUnolR+D
CiPEdFchkbk2oItnzf4Gg+DQ+wwK8fjrJot9fqRbzS4sba2519crOQx16FMNMCjw
S3giKzATd4iDKx4fCx9sLT3E9X3FIa9ezHAfsiLqPwkzeK0obn231eYvvQ09mexE
+fu50x+qvxV5T7n/H2EckTjx7sPr4+7TaIRvmzSAzRuoVOs/eR5CvDi4Mby2QpQX
tvw2Gs2S+uMjGcvWqF8prftV/QTuKEwivtbOK2/ERen9HizPQKC/HiH5Qbk0DO3Q
QegF6VztL4jHnbaY/uA+meQ/kMYxAnJIZjlGr1fRF0FMSC91h3spFbArwy+tvfVZ
3wnoqgGKfj5zIr5gkKPNgJpgJ3DPYBaAHuL7LnLx8sq+zkjX7UvizAgIBk1GDYPP
+h0H0BQZp7glhW7R9jKyS6iWIBWMq9rj1MyftSY9mlv06uDpkMrVR6hy7Gbh4tJg
8/b8tb6BXdvwppReF9jnK8BX6JMZgpMvZ7JGnzVaPq0TVsWVo6mp67+cFssRWXug
GkrQz43OqdCQ4wNOfGAXKV83j4nPknSmJ7R636ndnp1/ddw5ndSZ9pjbt64uZQo1
DqkoTUCnhyVtjvOSwf6DWf7dSMGuGTDKNb4TmEN5+eKn2y+Y0w9iscwKZ8GpS21l
Pfrq4Lipzia+7XgLLEzpwOwhI8fbZhKeO7qU39rkP1rQSAzEr3PDE7DbWxRq0SPi
jvgKtl/NUTGdTaQJsPQWf9+3KytAMEfoWTW4JOkwY3m5iWtNSy1ZiUcwMjHwU/Hl
xZWZ63DNPrGMtTorHwUxWhVwzndZbkIlUBLAyk2JF14LRbMH1ckeymjnQtNh144K
fsmW0Q9eSIkO/E+OkBx6xksYCwF2rfevSkJIc+VxeLWbMIpOSMueTO7acEORdIYc
Z3asxJkgAMUKsl5PweExEdPvZqf8aBi/ryB4PB63ApI7FQcxeHj2lSs/msT6KTnI
ge4mPguvXP7u5KuuchGVzeS+id5YMciwnwXbRttC2cKJyWtJYU6JKpbxtcxU7G3y
ti8AytPpgfRLVydWyupumrK7c2L+QA9oKS29njE09phBr3B+ANwzWa8MC0UjsVRw
eE52vTHLFb2iW4iI3Yu7QpHKQwDnn7LIonkZs3yo1MTINiXC7PJMxrAj6mI/Migm
HgwTsuhmRXxSFSmKpHd8YHsdj2K/hW+VzUWsGP/6vxGXW3TCk6jODN1JoFKdBYNd
MXFB5dMROi38Utr0AWDQDKOK9NQcGacfI5rZ18leWFUocC8wxcyQyVpI80OwcPC+
QfwTMXCdYY84plOU45oNpCZNXFneEMTHvTqeCr9kf3Y5ZMpqM6TYD8GbxT4RKPhi
RJ0/5nZ2gy3ZoUKn8OjJ21Kn3MUOrkqZRXlvi8vAdfMZlB/B7fRyDhojQmxzK4h/
ciGKggSqh7v2VhooFrstPJRQNxY0p6kPJp28OtZozqM7v2hLFLGOjYtD7OO9FCBK
svgkN3h20p/se51ETH3+GYymEIQjMzOdiSAEwyyTLcdfyNg0Mv23ZDugLwWefdlD
2CKWpp20NwkGUOqeRxqnYP5lEmu2E2XrVsJkRJHOh7/gi3gXeFtJ7o9kTxxgkXeI
jqoIxOCKWtw/NjIuONeeX5bSDPZDftFblRGbt/qHXdPhUjE5MNH9gJu3TOCyYJhd
WeNqB+Ku7R1PH1a3oggwy/Tx/zP6A/IwoYP1nReq23FlPhjscgfElAadZMDuG2cl
nFOG3z9KUGaPh0/ATmrsF/oE8QV7wt2HjpVv5ub3qjTLe7kALN2UJSwks18AFzi6
lqf7iRYHtdyuXdeL5rlW4qki4whIDxGCYXLnO8bnza4S0fPnEw79aB8B4oL9WkVD
VVO09mQLYtCpwwObYDBt8xV+rzlR28UuxREbKPwsqkNIMkbAC/L7Cud8kH7NV+NP
cBNKCS8Xz87NA9TzpixiOrBDzI0NP1AVcBk2qzapsHbZ3UzJqxoNBjvh47wixvAF
6SJrDnen2s/PTORJMIqGanFow2VfoDbQ/GXm0tgg51yVsBs0dfzY1+K2FIszcSnV
skFExG/z0n4ot9aOaqm05L1JOjiQVtjEiezuE6lZA5sGHkXQ3stEQQCawsIricX2
waIb6lDZAwljuoSm71Z1195HEyVzZ6gGpOdO2rRzvIE6HhdAkYCViYol9TG5R13K
y77mRixL5MlN/5ZEdB5GJ76rd8m4Yx0BBUYH8ozVQ7h6tJ3N6TFctvBpbxscFiD3
PsKR2XNyVw3eOn2nF9I/zwvqRg86dPgOSNIyQ9epelbczIsde5swzMfINVe2VVu9
M7B44BAkG7/IPO1PqfUdanW32yRO6BQ5J/OmnvE0QizQpHN8mzInoQnvWf231lHF
rTpPFUfaYmUGdGO01o8DlMQfi0V+m7VP4goz78tqRQ73sTErp+MsFn9X1vvfLoUI
EThM43fAsXYpTHmuwscXdCQSDwNtw+YLW049wVs7KoLE8sb4l+XxcZyGSVXcPFC1
zoF01EckovkRZabqsimkEXxpozwc1EOkGAaAsZPkVwPgboPajQoxfIVqBSETrdih
wWEm6yJrsKRM6zz2CyA++VQZL2S/Ayjauqjg5tL+gSrT4jmmU84O4bxu7PME9H8H
XRanT04rA69puNDOZkWBBxZ+F8ZYa/aZaRj2zvwSVAARj2slQvmRbjIemmgo09nM
1rZdi/dbOWcaITvpINvgDZewCvf1giF2VwDJNdR3gElxZF20who2XNozk50StyBv
yd1ZH/mzRUCm1qHrQ0DISOixsD4+klMXt3R4DU7WsdVhhjxTzWAhuya/zLZxlfZr
YpDO04/cr6cfBe8Gix+Qp6Km+miJhuYZu1ZwEDHhJ7SZ0/eS9zxytL3Ax2h93/cO
/pezz+r+LvwC8hwmY7IsSSYKGPBJ6TxK2nBlQphQiu7czvkp41/hOUuYUfyNqJLo
371+HA1QfpS6jk6YG/AoMuKRN9kD5AAGBWnOWoKfMzPECryFl8LmlBAZQb9rwP3x
LV6R3la8keXfbsV0iOtYP1eVbG/qt77Aw0Qb1Ju6Y6NtdEHjTMe2R5BCr9XznW8d
CbmFKL2+EGkH4Ib8aYdqBaT2QmI+hrqnfjg5QhbBhEr+GsgGfm7AYYFsVEIhHK04
yp+Hhf+Cd0uR0yHwHv/5uhGt7ePLTnTfC8sQQcKXPf3aoK3PVjtub4ffrNDdgswa
AVUZYhe2z1Pcjm+nw570u8OLEj85kpftzX6eH4VLtk2TtM77ziuGF2sFOeCgpw/W
te5qoE/VMOiaLeRLhd/sTMYLkhNH6YLWOZIg0q5hhL/wnt+zvzTzNAqd4eSjTaVQ
HNJL0gqwT6MunCAK7QS1bqVwleMB8jW/hAPQJmgC4S2GtlFbqeRngmvH0wP8v/4G
EnsRPcMBXYv4reXme1z1x0oCkjrH/IC+Z4t2LCIt0QkZrpbZjeOuPDuy35INL3L/
DpcTU6piY0kVJFSiwjaDNRFUj+Z1ipdqN9Hew+nBlf3HoaRBlHOvLKFYkpmJ5036
1kTWaDMmcx66D0msNhn0SgMPDNnzZGpv5EFrVdF9X6rfqgPQ2Ii+2SUcY89sxf73
I5coTY19p/9j/IEi1ToLqctxmufha3KTzalILWmerPCQQ8576NfD6nQqD35mRyNy
t2CLD0hpFbtdpCvTRd2MrJRusJW4aC23QHr2naGx0iPpz2VvG6lmAJvrZ7uB9Fz4
Y0cfhFuS6TXXcxZGdp8w6hLFpS2d77BwRWFUfYZp2vb+46L72DBovdJTeJ9AeACr
RcE0fbgcAVZbgVrl+q4SbppcE+Ud35/wOOohPcP1enLMMLLHGyEkvjNyww+VkfOi
VO0bF3Aqe/HNQi3BMYTzX/DVH+qi1uYzj9LEeJwQuwus9K7cFITmwiPWASXl7oza
IUmt4vh41fl404iT2ddQW+DSBjMVymegbU8jG51kPfsra8Oug+MMVVKQSQPgtCPn
dKWDK+SZuq1YiN2iaR8xWZ96vmaQwYHxEwgac4DXpuId3dT2gF/pHoLi71xuyLQ1
zotteBrhVshZ2FwOzNeOCHFLRDfxVE9/ffogme+NXvFxP9nGtR/FWQeYI/gsFZRY
F65ewedqAu2oAPh47uMkNx+AAZRSbq+UjTWXmmcHVMRjGMNkcu5CcBh0sDsr7MBB
7QesEfchLU9/j4LcJgUzSxJyoxj7W9lCHUSlns6fDSI5FtR7yhBitQOoEs8aK/3u
vmG+hXVUXyePRKBbFlVjTtq1cZbQy6ePQ36I1O8T6J2iPZ7WxHD2gjticumtba8p
hFqEq+R/sAK8JP6fFX2FVkh3dGQVQCd/Kufsta8tL7rd57AFyKqX0GRicFiVDucD
9/nHS8J4CW+aFKGMVfFAH6rIkfTDO9WYpc4rwUlKrWKAeEREPUjMZWj/Pvj33WSV
Gt53KmIfb5Rgb5SarWl0kg==
`protect END_PROTECTED
