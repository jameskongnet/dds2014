`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZR2O1mSDHVH2KA4OWgdSS+3WIY9n625fr5V4NWX/DUgrBGWI75O1IezSq4zC9frS
Q7HlQQw/uwrzpLD6RXTmoo226oYaO4Yau0rrsXaKIF6euHp4b/4QhYQB7eF/4erR
GwbpxaexpuqyZ8uAhgzvqH05KZLzuDBMZrehrtbDDXCdeY9GPCfVR8Ep8xvkGozR
dBtpCAvFzEZurGmZY1z2plbNxlzwyGLpEEXCb9/FKW2zQtgbO7sXY+illDDxsA2q
/YGa9zwDj0YwQ0UO1xlBJhS/l2758W3B68OaJegX7hSrDz0YWAFE3jpxKwC9vX1N
ES/FoPKdSReYkQ0BHeqnhi2QHx12UxbtNBnt9cbMSyB3O7oqkbdgOYlsiFcpLD2n
D3wa7Zele0XXxEnS+N3OM/cXvSb09HUtJbVB966rtru5TQtxap/3ktYWwM35PKm+
Tjc3xBy2kdAiZBfe07C2NDD4epDhn6ZX6PV5X+LeFAHoFxUs+aLUYYTve198XUbD
r86Du1cbk3tLT+V19d8RrGRV3xGOwHnOPH25d7lPIr3wpeiEUD7LKaQG63ttsxjL
UAepNS+Z4aBOc9AGMIFaIf0FI4P7ggx0dClHVRkxLDGxFYzvvjLAxp2I2ZGHNkOf
T1cghMXjdjB1KujAb5XH4fYSI72lx8PVUHzekc1/GWw=
`protect END_PROTECTED
