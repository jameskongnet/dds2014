`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6hRkSooeRrfpQ9DKBJAAexiDyf589+FJxKK+NDDkYMXj2OYFF/+Iwb3bZT15Mr0F
yH3ACi911XB29HLuksFBHwwIAKEOC9TbvphTmRmnJi1Xlvm+i8XAcs8ESvUhTfp2
bRxspJJjZ56Q2WutkODBR9vxMDVfLqQEyC44asehuq+Efmey0gOn3pj6Vg0uBq4I
/wXf4UoP6qX5A4WGmA/KNbnabiSg0JoPw2TuoIpLlhiholmbuxOUohBrOHTSPMNg
CC+n/Y/uHSJ0pyBt/5i+Y3VIFcpZgQuVywBa/To2wdYlg8HWAGOgusUXNeTwyTow
BYAtUWflT7oVaY4a7gQeSLZZICT3dkYBMJqCv8ZJIHm1M/8V47JfJlRO22FPKxiO
S225cJ8NaG3o/fwbHq4xi9rKSxOTWcSpfrNtZcqbmuu+FUx++l+IG3xdKG8JE6EM
wm9l1AugN++gXnJ/KBr/qFMfZ/LxC4nWYKfWa05av1pVqlL9hP77gvHkB5y9UTtq
EHKKl+PCE8xYQXgkrM8ol6mND3HebDWR4F5QvAhnClcAq8G4v2MmMr7KdC7xFojY
0bwJpjyqZzxkUrMK3c+hfE6b12Tr71foy80R0RFJbP1x92XAtt4WQSGho9uMsPuz
bM0679oE5zeb4RgCjtUNOil22p2M2mG0hHvbkunw2Mvu+0vB98x69coaHW6so+J/
m42dgo8SR5UxzSa2yxp4BrLMlVxqNc5COj5HkauZKMd/EdzlhXYVja950Ip5VqPP
wk2jb6zoFkwBj3CMThE3mqmkTlrktlrYVT1s5QYq47ppzo2wrqxpnPKtQGHZ1R0n
jRoJ46jwU2918qZ7OGNExNLXu4zuw66a7UCV033uhrlHqKGZB9yEbGeo99CckUqU
xJrELDqU9WabvqCo9MfykiYNYPABmeGUXVrCTXgJsalvyasQwBB1MIaHLKUZQxOY
dI9m1YV3in0APDIssa4srdKbxV650AmeyTPxYJHoRPX4t2ufnC5nGVrm3+kJbh5u
8ZaerHI+A+80g1W46jDm8zKck2yGryjxTeFBwMp60U55DFBG7HXJCpMavXDm/FAG
+mvuZHGYpL1rWpZ8FfQpeRsqleiUxyEObV4UixPEgdhnqoy0HjuKexm25k3n0n0e
L94Zgh7/g+/of56B1xHm2HFTdlH3NjGT0DPE8Ynr1DMaGMBkSjFPrYxnhIoyW4GT
s+w8wjc4b68i7lZCGQ3uePOvkBphFgaYvyRHr927TmUZDfh8QJk10/aYYLIlA8ja
/453/ixbFZfs33mmvT6W0bO9AhrGityp7XNMF49mmGwJBnbh0yYuPLGMIulP6bFr
f8JEv4BkDFIvSxAko3DdYxgy+e1fQWnMADgzk9jvSfEEwdDXWePzEkihYkWXAAAO
xCUYpadCCzBOnu6s5VzNXLFA/cyzFtvoxI1AmJctORZvAYDN23RjQFGEnwtFKiVE
a7Fi414XBItY2YH2AiK6+xZVd+LI3IeJ89gbIu9toX1FzJjdpgJG18iKVdrN3Oge
m6sBxIuO/fmSoVzJ9VSauteQNh+rsldVSxzfZV3Haa/0E+VAKblkQxYZQVuWB47K
htfG7+xn/QmCdmKicvkvzyBKikpszJ3KTCy7QnN43uk6r9aPpQT9Lyqb1YhTD/Y6
SSpZipxF+a8sfGtvJm7eQrb9BVYAGOOWewomjvaPhk5QldCsY8DpOiKO37h9kJtO
VnIgwtnPP8tSJ7/J4Ntuyz4oE85cYRkPwSVD0RNxY0nSDv+4D+xql852Ayss6ujO
zW/k+krPgBwwc8GR6kuYeO4JKcFi5P7NuQUT5AObpP/tF/ujxo6elPTVPGJ7/CSy
7F0u59AYcMg0CHUCe1UILs+k6uHdwR7c4KK1rMyowt7yH6cyy1nqJIjG4yNEbOzW
S7vFFCHdG2fx2IsznfEnCoDZvw0Gj9Gd+a3SvfNufbBGGWnE9QSHEz/Is3e5L7Cn
jKnZcycFy/+FE9C0ui8mU1bnv+y9ASn6qcUZTto3gr+p3YmaY1gLO8KEbefAE80N
IPmSNCxIyirTIu/WBQtbrB46aeLUIf9SKcgUMh6ki+MzqwUl1GR03SPb9YCATNZT
1tXkz369eHH5nhVPxoCBV2dZwhZ9Onpw/l+Yitxob9jI952I1H9w1S0zetiF4Qpx
aIFS/4cljRR2I2/spaKyrWlQWlWM0CJmc5lTYbDVVJ6QLUhDzupKxJowmSq6aAQ7
XCm2XUWu3Lk+mvRXGhAGNSAjLqaHP54SmWJltfNvMWGct0GVfoRZNAZ8hOtAYuEi
+jgCFH76u89//zV+yqeETIZjs7dHZkwf+rG+MhqQWqC9aGQoReCZ/41lhZt/XHKo
EDhF51bXj/NAQdREb2Q6UyMLmIwqe8R5A6PCg6O8mbJ63PyADAw6dvXx8Xa4yz89
CCpdJGQJXjMa5fE6AOLTpzI/+0H48u6jycbMBxF7HTfvwZXEWN1E3eGmEhWtI1EP
gvpoM+CixHGZDTHzfK+jzWo6ZX0tHdkgEMZdIxI4IikMssHrPP97LRR/zGxquZ4+
6b3KsVmO3fPzOSMuACT+3rXKByFZFR3NXRpoaM+xJxhps6geecKCLPvKw52nEyvl
g4Slm388kGkobcCP87hhrhFeRlnT+TUSuAcAdXQfPgVOcm7jmEh0VbD/h358HQl+
LmlGWY0fLoQTgvMi1su6CwueOSWdpVqbAvQj8Q71G3cZxhrXtWzKP5JGfBrrurcw
sAmFEa5fIMCZE2K4XqjOYWf9qS5WlO3Kze5yWHzphu3TiXAaLdYHyhCs6UNnpXyS
xGTpVkhsSDQ7ecNBYPO3saNadqV0Z3ZmO4x+rnEVmOQLr2OqS3o2hS90x5BSOAiw
ZgWbrDKK9Y4zvplFAX200S9ZiVaG9UiaahjRjMsfm9jQnioBt7h78EJGGnF4MKZ3
kbdQFJuKZJmMwCmQ9mC+6dInKoiqVfZoC1L/PW/ZyehNqdJhONzeHS9MfllmbRq0
BBTvzjDK54gtF1/ff7s/XpJ6pVnqvZ85bAnASYp99R3AOstbR/pbsm8seT4ots21
tA+7PTbm5Ecz7qmLEHHJYEer6SnRv5K/nBa093kCXcTMn9qqZi0OCVoqRdW466OG
S31SRrO7gGXoS5ABdebPnDMCpcS4UpFZGSD9uY7ko78MWS3piVpInc8xc55PbPPh
OTrQo5+/2pKatIBmn/IElyWJ9wMmS3OoGVe75PjSkf8y9mVEV6DpwPnuZ7PQmNAm
OOZGswR5ALqt/dwkWk9U385KbCKORleQ/4LMMA672Wy1ZA3lRBUHv3Sv7Bz3XIbq
fxSt5kHNDDJD16PK9Z5nKB5fmLVWHaOe9Dts0BQkRUUbXJnGi6smauPuntztJahE
`protect END_PROTECTED
