`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kk66YFFvmvSoJmQX+SBgCGSIR2yLlAMlYJIeXUTk88LmG7hJszqkUSi24U1XuzPn
7sihlc+rzkF9OvZDFnnPLIsvqus2aYzW3hGZl2tZhQKe338BBaYjKR5eauo48kVT
lSfhDVKECwsmWJeJCoQM8avcYriyevhRx66f2bKbbkYUcNwh1ivwMWBzh0mjFdfQ
YO73Zzmm40wH0SjnVjSdv6cFg5SrQ6BCi3Tk+iKNozMWT+Y31ulyIezNRW+KXVen
uAqQzhjrwlU+54HDkaPAc8jmiIkyJsI6EoJtHXdoRGeahGjJKQutCwbsNoM8eycK
wCZmZy/pxo5EZRLiCl4XP1fjnlBQBMOlSbP1lhRJFTpktTteYsOX8t60djWkKCMh
3trlRtOROjPIPY2wHM6eFdNoprdOxwDEF+mKf6eoT3OibKIQZ7n/IA/UaE9BaY4P
6nDLtj6w5TAy95VuYxLP/nRfU9lWdCNOySmNfvN65NDdW4QQv9bN9KRBmXtE1TmD
DyHgJgcsYTpKecK8Vo2kLWB2Bae5sksdFJaNHcWdKU84MibAp+Fr9+S4zG2QLRxf
ExSyuZHibe1FyNOI1davOM5ANWTyF7tOri7StGDeCt6tG8S0TvLTovICsD3KENM5
8xIz3zkXKywJyDIPcxrHNoPgLJj5YjuOO3HE0oLs9YsgoaKc3L80Gxl+5nMOHFWg
6rHRS6mnQvzREUYHvT/G05xFceyC5+4iw/iw9kHXQ5bEaerRZhwTTil57J7gsT0J
1dFxiSNJjwqlkfa7FKT20eZsSCmrBmYRvnPyJfnt6bjKCt7Y8QR9FXGVWdzZNV42
RjMR72BBSutP+oImNwDRU7x1HtjHfCCwGOsAF4BFHoh7YxFGl4lHD+u7rayd7d7G
zXRxRrkqV3QVtwmdHm//sLMQb9klLwuKTMUrRdC7rXw=
`protect END_PROTECTED
