`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EL02QeOdJJULAtwIj77bHgOcvAC665xpdw/fhip3LFUH+pN9+Tis1gJkLumYTVPq
3R7SvzrfpPV3GUQBUdXr1VI0VJU4L2/0TbeH5tvOBVcqiNRWis6UoHwFtGMeGxuI
HvGAlimRci6uDgBENjYygYQ9xkIKCXunDEPrtHSRw4ONBbkV/l+nL8YIth1TlGTa
OHizU4wPw9GnfG0+euJZrXhLcPJELNmHlaW7IbWCyZb/0mldJc0g28g7fLaloF93
C1txuMzdbrg9diXJXlAehGkHVHGFS1o48AxrRb7uakeoGcETUKBY7YeN+UcEbJEF
+le4HU21H+DnVyewnBVKRbSRJ7v8ns0U3sfeXvdI8Bc4g6brcPmN2TYb+78IIi/n
92S9vUIJROMYG5IunPUbR/jzyjmMF6nqTkqAIK9JJfC4BR4+nL4riiG1SJCIT9JE
WwG4lp3s65h5YHKWO3uUXE2K7zUzmEIvTBmN6jV1gnLXisDlWUpMcOCHhV/JEypR
cWKNJdeEdxjAFxsRRDEfDcukFrw+OhJpBabKCmIx62IKsqDv4dbZSvj1SY1jthA1
Y4YsCwWT0lwz2ulRSo+M6KxgtGNcngpb5Uk5i2tU6P6vlrxps7XdoEGJ5JHTwAcD
+aiUT/NuHQeanuQl4IK1iHkKcNFkPFqBQq13C0M7wnhnTvI35hwADcOWI0nT5WNg
zarqo6OXYbL9JZscamxJD+b9bp9wbj1Yc5mUYDpkKcxA79ikeRIKQ+8Ce9q38f1Q
ljKuDO7Y73cvboC1shv5kDJpFnuDapw7Dwu3C2U1V4Ar6kA3yy80nOQ3+9mYXWMj
WZBV+04Aau5AcM9gfSjSAuDUVbilU6EMBOc7HL20SMUm0etl+9QG0jqBf9p+AWB6
FI1nO8Zwum+f82co0cCvkyHMoGIIN0a8SItVvShP+Eui+2NGBSoDDc6wSUvDje/F
YQ1O/dTj7IGIT3M3zG/Zf8hrF55X5dq02beGvrVcGyTefmjNK4/8h8Qtp1gZsl5j
1xQ4xoKsxI70N8h1t8lLJzy+nY68lsEIdnKOXS0v5klxu9QF2YtLdzHB0VQIt1yR
T7fNjZr3KnvcF3M1PiKjq4kPsTwDlkmMOqLK/1ge5/4AKxxwugWNZaCg6zKvIbcC
He8s8esH/pBrhlGxYkUHAjw5UvRworIwzNDdAUbp2qPvhcAEmk+j7IfWzff8LL3V
rnvkwpAvcMQ9Z45Ao2GjtxJNO4SrOgjyoVBBtAz36rUCaLuFWnqtx1jFpN9vRszQ
5x/VbEzU8wCT92HHW0vblwANB/AiVrmI5pGLEabIJg5WFXRMl/XqvHTg30TOdHpg
pX9p6Ztd9YwVyJE7Y/d372q/40vY2f72Rd+ehSFu6J4ywgJFNdI+v03Gt3anUGb2
GJizdH89daxV+F06r1BjCgBJCdYnWWTr1i8K6tg2HNveBJWCYVS/sILmR4Ck2iNT
yKACB10yU/SZCNNY26YrtiMqxh+KQd47iaGvv0Uzg/QyIir7Vo5+aO46MxcSOc/u
iasSQnh9xJ1Pk5wPCVbVu4As1ZdRncgaOygQ5h22KC+R5TUfVN1cw3I5lgyCxRwA
44dIdGC13qnzD6dPdztHvv+EY6xn3ye3KL4lj1yuW/r5qPZJ+CkQilenXZz4TZag
WyQrZfMGYJCmUmNgxctVCwW4dc8aX0VEC/0UWMrnHdGUWQROD9h/agGI2VOryq1z
RrfHlcBkThYyZ8VBuN5kYqrtoVj01JTIYYJthPbwjUr5H0j1KzpS6cbPkyHSkahM
/WnxaX4whzi3HywKqq7wDjrZf6wEYF+eSI1kKO/fAvur3P3XahlFNwpwx/0e25Oe
KT20uv1KliQhru56NR+fDLoUv2EIuPhWkJRbUrpcDmnZAcki683s4dyJjHitDHp8
QWv1dtEWJHC9zAiw5U9QXpVpeDFICRTzyyVXlRsHlWtAwYebEJGz4tzDoYfncVz7
6T9IfLRQK6JRrElmwQeqnbs6wfnU33iKFxRWDNNMWTcwKcIYGt378Bk/n3Bjfz4T
PbhiYtlba8ZKBbFHIfZsogA66O7IoW3yd4VIxrFMdSnpYJw5wGcuVUDiTXYjxKnV
RWmROKUAGIrnsgSZq8XWbCBqfRPCOhVBF2x5ZfnYC/Tlo0EBKNGRZA3giNLwFBPv
2bALRjfGPpgOQb0J3Q+lvu8Y0wuDfEhXr7cojW4srQyfFiRn/bWiSZTnmQZxW2Co
VR+0TSCM+RKAoy0Vd3hRyQWIg3ghEwvk6/Q2a2yf3U4D+fAT36EDx62yA+uLILNu
4F05TjYB/d7q4wPIZvuGvBPMCgXXrxFi50HlAhfUkw0HhaPhnWZggGcvClgy0BVI
yygQ8dNp19kB06B2s5tgaP+rw6wqWj1yoA+ucELJXBzrPTIl0+WiynWnHf9HJxOJ
U/thEN0SCq7jBjGYK288QIexAVYPyIsxCQ6D9pny5rLLZbH4aVjJI1+hlUKRCXYU
bdjEdcaAJNLoMZq6JzJOgguxE6hEYSTKkO6UPIaO5HGXNNpRAj11Mtrc0saWTWE2
6K0YxIl1OLjvSYvfjXjckL1fKAdt/whkdiQSuonturyRWl9ufvQwYDdhgfrHVWBP
PnPCyvbbtRTPZi9cYh29SFxI3Mo2BuwK9ZCGZGVh12j20diLV4+WWCSa82oPZLYN
o2USY6maBtNDuyEZIWnDZDn1iBR6LHUzevGTpOBXS8LJe1El4EXjqIvPOwsWFwQ6
gXVPSrT5fu2fMncP05zRZkqK5Eb7UG7CZMLbj7dqhu+C0h5/sQX5F7BHVv9/kXLt
H3SLh3L7cEWBdlC23z94Q7VrBxNzbB1OYL3vdKu35+/5mvrO76ffNiaU8SZq18F+
xk29dIvcozK9qpW4r2MOKkcJ6iI5EEAEbSbLrM4VAXrJkCLX22j0PbO2Iovm1xow
m4yARD+oM9+pVphR+tW89o6efpLY+0A02Hfh1NZPUrA36EWQ2lPcUhHL2S1uWlna
fkRqfRpTAwF4Lfr7xfzpveyiM4sgsY4rtGS9ArhU0OMW0q6BZwSnBGrd2D/LY35g
VEjuMOEG0xWmvPecAcXrLAuR7xQB/6GvOwoOS5vyX7To9Gt3FOwJ83Cz8vjNHo52
mZzwdUgtfODBw6pGK47IhN34jEB9SoHVjb0gbq5OUM/M4syXK9MStBixYce/j4pW
9SOiLzWb7TVo340NtD2uRl7TicoyzCPt/CMHbGbCcphfZsgR3tDOGwi/GlmPaUnP
xhpqoOtE3TKqodBK8m38FLurFbUFHJmIG6Cxktpy0GH2ieG3vI9RV4i8w0ipnnSo
uHx0PsDTkrkiAQIgyEiUn/LSv9jvWlMqdCmBJChdF5XhfL5tdHF6aizvN1E7AWh3
PmSR6JN7SsDd5X01djdlg5+TJLkUAP5lSxfsoogCi5zUtPYNlSo/r+YT2nvxHR76
xiL6gY+OG1Ekbi3vTJzrYCerSFlcTztH8ENQXhnsNcr1QI7XPAWTRnXJFaAw2+CD
KURdtqtCRY6BEMWSMXG56mgYioqW/o7ssC9kXjLSyI6LFR5hEFEN1GOnLLc4h16g
BaTl4+QqQLYW7pGuNPb6yFiEyqle9ycrEstO3IJ0Raak3aXrFwHTRqrtZfDLoxNz
8wgD/PtiKnna70VHhySzfp03AyYay+yAz6wc+iYgKJrCk+5RCWTUFbXaW18C8ZWh
L45EBNd0ptiAWGYSkTvk9zaBJJoEZe/XYRs6c6CiEa9HM0zSHj3mOPUBnBX9yJe/
Kqq6w0WRfjo6IN6Zg360fMIHDTwRqmjnrpDA/CfwHFFLHMTvWDQ1soqfHmlEQBfW
Lt/I/bXXYWZXKjNscZ+YrhihYbPtkpnjwZ2qsO3m+bz9aHB37ZZ8qQqoYwHqHkOe
zrGEntOYygkS8Evyu6bJ1PkL/MCIa4855pydOOUjiJXWTheCsTM6uBUX3EOv12+O
76bLxdd8l1znkI8dmxl5JDNVd27mPCleyxtPGraJhIeXTqGSXUNjWNjNzra3DYBQ
+HibHgo+90Q2GGrdQcx0HvSEm3LkGe1vxW8LPp3vtOIhR/fAzQO8EXmF52jaSMW7
Eq8pomet+43K4Y0RX8e9v+lLSQS6cswJ+1rWg/yRFUV477ddeR9mtApFpqInJWAf
lUlYqUCLQ9Oi1Mgxxmws+ocC9FtmUXw3kA9ORw+pernrf70ZQ+j/9Idc4JFlLzyP
fMjexGs6Y0K5zBcp4QuEX2xwUxF2Yz8NocNIXDGlOT2UlLHWuheGHHPLFbyMVZLM
Sp6dsTn5kyvn4ySM/uU2BIevtXtjKf/lC9gDOeSLyCHsxHHiBQ13k4aLCumcJyuZ
xi63YG2cM4LaKFFhCJKg/U0A6ZrGWxGlAfuGi9ye2uBIEhYgCVIPqxBjL6nCb8Qa
+GbNJHoQD11ioQ2on30cJtA/H+Z3GnX5PtqY2F1aQ67VlDEhd5+sBVes5NCCWlxr
C2BGCHztf/n21v6QpcpcmPxKw4wa1qURFWD9dT7yJHtSpfrL6mNh8/qLSSjBQfII
sG1lqKD611HtpV343Zi4VcsOpHqR7N9kPfw8e5Ph1+kIyJaXqfVBM3xVtzH+2V3K
wm8QMmyicw/wPoRO7xGWmS6JI+0Kk/NlcsQExLz98eCtNtj6jWB8oW9rx0oEVIja
FwFIqx77Y50LnhkYtloD+bqWVExE/EDKZouYoSbiO/xMTTw02sxgLhgTKXf7Xq8u
lam5r8IpsMkrsVTh7AnpZi7H3SbH6RZgm9VhEEXxk8YNU/dLQuRatTY7NWucgkYo
ne/2Y/GvpgPIhgCxFlYBKfO4FfKXWamJR4xC9DCBW5Nc7Uj8Z9pEB/XaOBXimGLY
fneBiI+qX1aTbMJwhx3YkzkNIj6Km+kf9MIZn8QJX/b3xKeyar6vwXepbJX4Ip6H
/KGvPS/pOsmy8U6VCcfPeqf7h7L1/rAAKHjEqqONMv1jr57SS9ckWLqUD0m8qOfN
XGp9JpNMvIunlf0Dc4u2t9fDK+zPwVb5AM1wSEjXkDJ3kbrJT3R/ryrtZXSfUv86
dET3XgR72pTjp8udYbtmX2K5yPJBltMHNw/Rlb3bj/BCd6fEirZqDxrEnKs3LsUA
X6Jr6R0+7xYqunC04bGrJM4Nb28XwY2ADH88nIGFtmJxYvgJTDUwUyMi+dmlyzB9
PK/s2YwEXPVzZrpFDfG1MuonkUT4WjzlxiilXHDZHu3bs0HEqxIQzH7LU6NRS4jU
99la+l2pxc+MWv5z9BU5dhKJFHB+ICMZpt++NegzPbzxqy7oZAeZZImGezIAG9W4
zekenGibOZgujUzqeiyCr2yYotMEgRHVeQ7Q2VBMIFgmxwyt76TpezHx/q94vv6s
9GXQF/qSX1CgG/cd8c2ak1rFKPw0RXijP+w0VXFF0GWN4rJ9YPkpjaoXVyhazaRI
SrEBNoHeEBx6LJamOl1mWakAZ9Zv2T7UQKT6OWX87+zGmnkqGZeLg4yXHkAjRG+u
MMiJ1PokD6xfzbg4go84p8qGDQ+mo7PKhy3cktMW3mbSEJbeQ2V3cW2hbENoqAwh
oGc28T0la/szpmeE8BUm4rLGRudmSFOaRVtndEpI+mIZGXN/1v88Ye8umNwReyOb
QS6JqrhgaZ5Ancu3iXYKdjhdVMR0Ifv5lJl01h7Red8IU4tJFN8QPhEiitgIARy2
QqPf62+mjXLifRs774SkLPGL8o2GnA9EKh5pa+g4iOpgWlKJD9nxhjXAczeDHLe1
hWGIy6FAYM/0MczZpsCaoC4qJUymG4NwXfZIwWaMGmcq9wU9xNL0Ix/VxvzC2n0n
XAi1fEcA45kJGrBVtIUBZ1TjNwigY/FvmCMPl4dX3MdfxafJmpHTJQnGrBfyJ4iy
eU8sfEB91/bl6xh/mwCapYnbHYF9CMZgo7/Wyh3Y4U26EOAaFaxTpls2b5mpSEvO
oap9CyT5mp6PcaRE7dXh1FjNkt7itettbCMARgmXSizmNwNRi0i38lpQAyGHVA/9
S12Kx+H3Fy3LAe9XyfjOMpeDhDwVHkmYJ9T3jvuSuP3t1h1cX9vDJo8X/fNAfPEx
DVxXwRArhKnp3frVKL1CyeQljbFuGJ+1ixhOQDTToW6PEah8lmnxX2j5TigAjlMb
HHl0BnDnW0wgfcUlFNBozrF45MQN6XBy1mjZyWpMUfdZq7oOefLI1zupp/O9JA4P
YXMbLmIaO6zK9KibGIjBqYL3LDxguJDUkhuUjGpt/IOC/59nhNuEbND8Vf2DBpDt
Pxox32XSAYGQbcddXDiEF0ZvCUSEhLPX1ZCJtosMw1xxIfopyOppHeQoETpeFQ4o
7+gy6jh46GQP6Z4PPtCiaORWzS3kxcdpDnIo6pAEuoMwecAYRgFpt3QGyT5s17Hq
icfjB1umyuUa+2GMVy7No+j6efzjX5miZajt8A8eb54puJG62kDYlvfpHmZBuzIG
Yuk/jr/2hRGtM+MdUgumu/g7VHI2DmTpj5+/UstG4XtDaIcImBT5uaj0m+zv+Ys1
XHEzZe5hedb6Ow6kDEacnWlpVT9EKjg4saB2Dnnxwdi9muLS+PkmduIByA/iu3/6
o54wcZgBsyhYAvqFf0WLJRPi0icQlT6E4A4fdSF7bfHr48YSXl4LuqnZ4cySF7iN
LMd1GcR1yC4AtAbdsmfIdWbxpAd2qTF6zpMupWGzdIXy7XWc7I5nA2OSEcq5oT4l
Pq8w55K6ssIYdTWqOK6R2Ug2/hnwDB+tmQHaTdxF7NLdA3skBjEiHzXG8N52N5yA
2qEiaEugrcazlGC4ufDxme0d3ZIM50diSaR+YmCC4jDZsvoFN7n5+plz9DeCReL4
YpKbawN8xC+vqC8RFJEhs0On/EVOly4DEi6UGmGhakcC6Wc5nLXEHe620qvP18Hg
AdaAT6MC3VKCNjolMgbd4ylWkD4zZ49Xb9w3mtyYpOHAPNH6YZXOn+Lu3RWjgzeH
aNx6TMABWhaGaRvg2fXfqLK4CCglxDVARRh33Fz2s9qvj9HM61N+Vwe2o8HUu/h1
Js/bzgjgIR/VqbK5U8wPjhw7hmYFcbRdDuMZFB8INLhOeLa9siuK+zZcNO0aT9Ah
nOQXMb5tWNw2Nyih6ySDrKxByoQHAhy6ZqaLV5i3wllnHVthbcJQ4mMYTTEcbTnV
CbG+skIfbqKHmwsogzCk3kB1kD8HzZ1bJuOApNOsaWoVxg8F5Wd4SmZE+b/K5/AJ
Btt5KcuH91mR6KB7eunxSdlni7JDM7qeB+tkBeg7csf4T0oTTwVr6UBxLuwOcws1
yvuhIRx5fvfivznpANFjvAQM7XUT8iPi3KXOUvTq6/PPv/tAQCjPQQCzqxKKWhEs
ZsuV6F8vKN0O8vipUGQIgIht/4IsuIXaEtLSW6RTIRtOIegJIDuxJIEyYENzvlQG
83XpRLTT7NlTwjgB7+TagQ2wE2K6YjjUA2UVLxiJDX3P/kmiYIQbbBDSMwFSGU+A
sOLzuFj7wHKFna0CKffRwMOP0kJAG4tb69i1yqNUnMy6eAsvorTSNPB8fxQjQkEC
uTC32tGhWxAU4X+6wHpBAuBu898UoeqNKeOFLLQ9xUD0XKB6NZIIc0/xJTgJAUMv
HWSsQfg6dMKwUqstYN3OCIoGlhEdL6gIX9XIfdOJpAvWc7tNh7MoOUa8Yd3vfqxj
jUpZMbH/jYNi+CcZ3ghRwpaeXGNxTRkroatkowtDaKzJ/Euxpeiz8D0+OGaGo7ny
hmSxG3l79QQcFGyEv6FNgDPbC0N/OHMmSKrIdZlTRhW2gzOgWSFt1/3eOEHLSYJ8
B1VjOi6798mWAHKN3JoxyZy2dYm2U7rHm/05dHlyja3qvoJo6yLF08Im9UMsmS9Q
cLN6LU40p3md03tooCfKXDdSzG+VV8XND3V/F8Lq9mqpOEDMTMHyypMqoO4yyWt7
1me+UinVv2wxxNSFVHLukJp6H2lv/mFo/B1tjOuW7O89btz341cBc1cSKPsDmnir
P61sjWzMCVr1YiI/8pWYO5LzrVK+X+vRD7ragLIJSlIhy44SEufqoJqT3Nzrwkun
lViCTyU2veNPnOwXMS96lgxZe9Zhuj9xB+w+QqBrNa1iSd2V7JVcYgWGQLz2XQyV
HppblwOWXuVvcNKt0ayT4gXvm72amHmNuK9ej2wtOYWq6z41jWxKsAY8xSBF1hYq
f6dOnR2qHgxKPrcjifqjTrP7bBfb7/kODtXSJQTqfHMcRbeZmJJGN4W73mt3dfEn
SC4Z8cPB3FyTD2T52RxdevamXDLnkyJy1rktS8kevZkQvS/3G5n8z/BGZqih0TDK
Bc7T3icCXkqRnYApZgMVr3JUYPKC4fe78rn8qDamplg7EX99uEp0FSYbZFioD0t6
Zr2Oac1OB80P5CflRY31Fn2RD6JtfkEaF2lShW6FZLI0p+RcPcVVrc5p9LNQpw4m
OQDrvohPnV/sHymH3VtQntYppYWPmOC+dbxmG+dyXyVwIJgQ9PQZIWl40XU2O999
Qnv72r3YKtxC5oTa2RCoP/nlU6mrL2BEmJBEstE27MzCJbElXdfNVv9JstrdJ86E
p8gjXtfdVRa0lBHSGI5wYxI3JhqftGLYvJjgpnCPE8ydEm3VQeLY95+fJegIUD+D
qAWqyeUk9y4eY/60KhmjbPQYHhoyRBG1H8cIInPOm09DkrBKWnXawr473d9hpmPb
WFtMljxFeyNVHTIypOo1bwjBgF+qyj84jpij+OWX34jsMZNi9mhMdI3lavcVMPJr
rJYS1C5tX9GVkfMBwKN42gSCwOJnflaphNxp54wWsXy5h0cqKqlW8gxHoDzlCHFo
vy594h/xAc0wIsdQznuFQCrepTwr86j6l87Yacaj5hb0NmnB3VB+PBGuKhaDNEfZ
8jjxXUo+yiaf44jQSpOMNn7U5ff/tlBKS0QBtm+aSF015miqRbxlace4aFacRY33
smDBZbX2p+Ivvld5bJdN6Dc9a0R/IPW0VIn+M6zUpgyPMs5oLieb9eeP/2q9QwCb
NMT63Wug6MS0bip050W1/fRyy+2TdNkRGCoiupECf9pXm8/q52d8d4NI6sY9g0WI
J6mDBI5FcxuVUOXYL6I41v/fCLYC4Ih/faMWVpvDsRXw4vKRs8qK1/AbLyCoTSQQ
fOJyDzLSK3Lah81OVw4L3UmqGZZPNAi3fswDR99AWzSnddLjNFhak7I85XDPetuq
eQn1esYVVRf3rmow+rJHr/bRffokfFZ0LsZwymYNHqa4jAbBDXLJ9HZ+emJ+3C3g
CTqHsF/kq36ikT9CWrfibmTIx3gRfwXGR3fME8vnBBsulPQDUcgecAKJcG9EfjH6
dz5G6JxbJJrBW66NQcYbX+f7dDuY+msQ5z3CdVB2ReE6lnwfdoYPNlXdFN0t3ogn
wFD91oLF2XqJlFDA575PGJ/YVUGMlP8XHVc8mk2ZT3avIt53Gb381q8q3G74BPTW
SQWLi9uSRieBIuSncC/ss3kNtBimjOpGAGKk9y4PWRsMOf/er/YLh5mu2p8Cbxwi
8D76vFL67B6ourT9bg1s+NN2hPRhTArx5xMYwskIr0vEQz5KmG2OfM56EAqELIaG
DOBtLJXHzPxM7LV6Ww3LBoTjHQvoMRkszInl6xXy5DPHJpr6ulV0xmv2w+mOZARU
ZC3i3dPmEE1HZ/c5avjVv7gEnphrBtlBa5VK1owj0WlvDJq4iWCRTIZgjBU5Eb78
oJT8lROQuTwiPM0nrwvhlrWp9bydVfZaCUbfgZdQCZyyltiqoV5wg7hjwBX5kPr/
eHmt4jktdRNrMgZl8Od0PwVCK0NoiOruch+G69km6Pk5d9GuXBW3rNS4BWbl37Kq
GLWKCF30qyKJvvAewuw2N1LaiSunzubMfIQ1jNHMKvufINAS4RdCLNlLbWbSBNC+
OYZQmsh5Fqnmu1M2LWM1AnuuTQO6WbrpDMnngQLTLOfkvho3Cgv8YPV0RktBb8SD
0c8dz+vrSepTc1IUXMDeloosoxg5XyFbzZc8H896QmYF4uzcR4XyesymzdI8mHLv
7RLz2zrTZ40wX48HU6mc43RoroCeJs64XOJ1tqGd/Uz/fTZtBSg5HqQQrTVOu5fH
7gfaEPDKMf2p1YvumwDVKdntMRuf1LU5HwQH4RC7Y3A5KcbfObk6/w8sjuJ7dMPj
aEdnYVDrojQ9b9tGdCwWElwLOJchcYULzQE0rvR8kWEPh0eJToN5ZYRY1/ai+jWC
ovzGeB5nvHWExqJ+qDHlnxwumYUXDHjB6TRyE/mY1z0pnI7NvCY/JYR8AZhe2sn2
XkdUUd0GlL8b7t5kQzgVcVQ4cWeWtNBuvVGiwJk4gbN4erE7KLZfKWDpBIiqqo23
i1155WeFb4fGyc2rh4EZyMU8VWfmFVXqWevKte19JJPVBfvk8T0k+M76Sty5pafA
VEy/7XSJhKrIidM6E6FxJPuKpS5COqGBY1Euep9u/xap7F2ki1zSAdu9wmomcGUM
urISiTnE1MHYP6DUJKa2d81TIwEi50T78Kuz+VQ1v2IvHVWyp5WQ6+KPoaNaDXwq
ZTnu9NFmKwfn/UTftJaoWZNw1xw6ISi1w0ZHKvPFMyMMctjQwxDfAzcIjlbbt29g
OGmLZSn5BXXCNo/nb11Gwr9J8oMeXym2gfin9eICL+BrgyU9Jp/eBYitYACRWrJv
9EGG81CFfK6MhvqpG5fCPVHOiazXKotwe/0qFKRrvg4rnc1m1RcbSYoSJen2YlYG
mLmRIsT3I+TYcMNpRRYB5hfEFzygdDMMJNb1lRNC6hP0OTrqrsOfKaEzPQZ35PgM
7lbMkM38f1xDTFdqf/iapkzLPOxknNg1dH2YzC5NgWGJAUmsE0VXP9ZMxjqz/J8W
HFrzJ1xgk0fvAeftde6LRmt2wRCas8QyMBEO/DTRcOsWAbWrDD+t7ELE32fSOrrB
Z5SYK7xqSIIFYOt8ZswZqAr5iqAFmmEh/gmD39MxnTwqSlTwckXxjh+MzICPjhPv
RPPvoHRvrGViBBsIkZov3g/nl/dBJJ5AgY7yFt6ZnutY/KZSMdjbaJ4/mJH1Dox4
RNHZQ6feBqCnh6ZnR4b7S6ue882DZ0v6TAfZJmeetOvuxu6Q5dVDZ3MswnFNLBi5
uYInbBFUtG/gn7LM9K1FUbZ51AejCfatFIRvy3uHrt8SaZj7LMM+KRn/j5aZU3fI
Xx3dWbBIERvgcVOs5hRCa0gI4skrfN+z7RqC/jGSBl6+1fAAMhBUQ6mQXoOI1QiS
l9BNKZ4yt7EHGSAiS8LEPQReoJ+IUnzxGjewAHBAcNZ1r3zeWxheCYxKf5RWIzYX
WuPQeYVTC0pN89Utmw8JV4LHv/rKkIR/ePgx1qM+um+8VD0mSs+XRHjp4qfkFif3
RAKg5lLWt+dSTb4BaVy2myo7hXk+Gj7HjXMyCX9vkhKzANURHe8Cx6Xdb34oEMoH
Yqodto5bHmR1WGggwZzyHXmjM2VEAv7MmM43qAdNRXFDdAnMpEi6ptf0JTHf3gah
XXokJ8OdSC5HzTKpvdl/l6NXYMHFuLHEcWu+K6pQNkgpb/YGqtiScKxuFYJJTomV
QEzhQlDOXcEDvqa0ExpQihFTNg3cNbjQ6DIy3/5wQqLpdcwz30q1nSgBQKReoaF/
WvI2b8riksSdZO8RZgCNzXNf5pyBWqC0rsWpFyCeslx1j78SvbGV5PMNuMuLtxlU
T+5AtMHIvvYvIgwRTU4gHM/KLEMoTUK51V3MQJLXGMX3bF3YYI6H1x7DbAXDiSWZ
QnHk2tmkaqZ7gIDX+OKPm5/+wdTGM/nP5lZ14CPt2SmKtSruuNZgWGUy9jaQNKs/
lu7rcU4ok/tXstrWnG1/NZRhiUNsZw7HQiTcYHuTx0pN5B5JES8/zReLvxbVhigM
itB6/e6oNTBoTBsQulDX3LTpJziREjQqcTQo2gl5x/nXdRQkA+a2EIxbc/AvMA5f
uEFcd6cvhoms4jAZ0KNwhM2Ys0SxuoSvyXkDMdV4gRVHUfWbbu7NgpXT1k8NUK8d
7lFrf1Lv8r+4PnaOn3T1aQMGSL7CQ3ZZYGlgabc9bauVgYY7SgY4z8ThWTmivoh3
d5FxgkQo4eNg7ZcG4DtpJzcffWAhhWRopciLCkkAxuVdlhYIHl/rV1z/Z+i63Wqs
S86SgUVbozPN+g9PJ6BeLfgqLtk2dmqZhRYoy9TDtnx5Myo19GUbonWJCMV1CC+3
um51wmV2Y1bTfRrbT5IS80/15SRTpnZvZkfqULvC6LoFrNbOcp6sgk3j/w1HW97a
+N2uoqYKuTDjAtMsTGwcUH3VixyAdLmwS8I0EPQ9fdRR9TwRHeDxWDXo+qM3OD8u
puR2DmDt0iy1wMydiG1ysKDy9Hzic8e8j/2CtD9GfK3DKl+jGN4mmj2HYF1pYg8w
sKVHx1rs1MafyWZKq9vO4h/jKIBpfZDK74wU+4RmSkrdQd1bu5R4BNOQ2kwINvM9
jGkZFRtVR6JBa8fFQ+mZ+kU+bKYuiTzi5PATQxhRFLbIvuqYzEtFRC4mIovqRhFv
jQ9GiTkGjg2TBAnOoBIeIwlVhINyob+bu9C1ajCWAtVfrlLcv6a+0EZc8wyCGW5u
qKVMIfDtL9GZSfViwO3KBfIWOCGg9oCFPA/d0E0LDAmrWtTL50xkuyut+PYHDuCK
ZLcY6i7DqdG07m/5/Rr0a30txpFg+aRn59MtvXMwkK2F/jGyk658bC5pMpAon3Az
HF/eHmlm+oIN2C/Om7td5mnNCJQMIfj7CppiFXqtdQuD2Rn6mZ724hulC+t+OAWg
3vGEufxhzAtjgZno7vSW8GV1SiJLift1CIoXOaUbwt0l3G+Yr5IQtt1EH2D8wmj9
Kzt9JsddccQYjzAbE3/q28LRf9QccA/uFwOIcT0xNa7+di6gCA47+Y68D92vuP0H
/tPflV4AZE0eeuEpD/zIx91uElb12zYamMDxHk0ygO/ammknyrVmspvE5F1c2wdA
QqF0LhzPcyMdGutwziFVAyjBJQJh+mu4R5utvwcO/AYYwLcWNHzfKZs74eAp63yg
zfkUL/hejQoPAc51QQoRIPnevp75NXQE0uO8da3VAt91qXJr8SRwjkAHMBnJqd9E
NHM+0XP9SXdxOaGpTlGVdQr6dTgeaxg3vqNw3+52+QJRew6pJ9eXN+M4P6p99J7a
6IdmItRcfZo9XJ2pkSrNJq2et4gyf5WNv0Rg9HhlwtV1BDljy1JUNyH1XmRi6MPS
+YNBYq3WdbPincZAjwLmt+zdwd7X17zPWUhix3edGgxRC2fu/CXdbe2Zpus8wNQv
OAK+prE6TPodSVNdfvdgjw2PnH3d1q18MSMN+ydqDl2XHmTInyR10yHey+xtkzhb
wyIrRNp22eqxwxahfdeHWAgEXofLzSqbvZco+vka4TYUPS7u7qhSzOEn62SPQ5cC
HCqOfVZSOyou0NnAZ/6Au7sTs+Gyce+7gAuhAg5qA0k8fX+XosKB9GAPaEshNYHu
dX7B9lbd2NZkovkWkccxuFQhBSwZflk5RHO9Qzxfia/EXLycC6CKl1/m8idEk1l0
epm/aFkbqWBSpHyxpr2c9ahDqHpasiWOBFkblqjZn74iUwBGkoNtm+f2gvHHoEb+
FqRi4Y1f6iBdiZY8KgX50/SauYF1hAiLr8DJnu4H2jlgHw5TlK6kjQ07nGJy31q+
ZbFNuxkB+/kArWgeOt28VAl07ewruW11LfYCtUI4IkTaQ/iN317J1eCZ9uyYaSzE
vWa38u3jkVhLSMc0lGs1Lu84ZHRh8YADx0rXT8BH55A9UaIRs5O2FRmjd/mNHKC0
Y3pQhMaPDFCD/Zu6ZYFgCOxgETbvAcBHCgDfmz0czmH1uqDewGiVQsRXhqtyFXjj
r30xAUi060nyc6hXUemM2DROkWbqJ2S/U4iEkpC1lZy9buYm9p6ufHAR4Xfynf+y
pIGnXjVJJHmGLMV6KIEPJOXzUMn9KeK4mQSoa0g45TbEhRqZkM/8AnGqbs99Aigv
SKLu5LWhzUpa2n7UGwnVofynck7pIonk7M4QQWqUxU9Hv7EHB6yZ7R8H3uuYygKM
MiaraUecsbKQhC9SB8o1ax9OhX5U6SCqig64zk5HK5NawNYBbxMtiF1FTZJ788HK
Sf76L4Wkg/szixPtIb7lwAbgwxZ1TH4PhErt0Hn0yJJ/DTZDUFS4tSFZdpGGUsaU
GziSK55ttxQKGgqiVrvG+2b6NOoJkdf34mXvWTDxvnum+UWDlzExNGTv4FliW4xc
M8VunOcmXPjP0G6k/N3HaCQx/5khFu6E5/Z9WLBHhk4fZ0L1OxnLeZYqEmPfDn1a
5ZVkTsBRsCxAxrXVt+R5T2BceP00GP9QCcXPseBuELEow5/Fmj+lFjdZBLE+lkUw
QIrSOAB2tn+n2a2jmt2u/JxaKNZKmDmIn9ZtXmf6hERHzIvTNYW9aM8mAPXPrT1F
FCo8bOIHsvTS29GAOcrHiH0EU+w4KlnQowwhSmd5Ntf+h58hD0AyxwYzItiffd3L
i7TBHhZPD9f4TOE6wfykr+ICDfga6OQC9VCPBsSFntNNQ2CDcc8rQfBgc9BnjNnZ
gOOs4qAAgvs36lNiNxFsZRQ1+WsOCRfJwcFqi5pUejaTm5r+CZgavUSoennUdNX5
bU2wy7CYsf6BOfok+d5wJGdiB5vVOvUUllH/9E8d2YOaC7SEbhbSYb6mHq6CzvRX
kYzEaXDVAixWdSELnwZJ6Q==
`protect END_PROTECTED
