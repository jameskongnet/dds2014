`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWeqTxAKt9Ifr8wACIVXUGKjYmFIY18rnBiTB8OZ/9e05vsnw/Yv7pV2uMUBVibI
D3618weYbqOYP4yGPMsuklBvNn9Z8D1NN9SdP6jDZAr8KZ/1YeSxpJA8xaSmVElb
3zBof/rciot5YzeLAYHyqiHJKqAmo1Y7Y06YOBiJ7/PtA0nbfv9Y3vBNExCbaUqP
O1je445k5aM8igUVXAfnEWxcXYDXKba9tbr9NAE3OTeWgRs9MHT37QxlVzrUr2fc
ChUfw4yrWqQvF7s3q0a9gTi9ocIb1PnD+3v4kPrGyD4sZOlWXN/zLfsCqi3Voqau
tbdSERCeLNC6mWodw2cuw6BRGQCFp7gL18Jei6F1PitAffk7+Egm6++flMeczUR6
+Ll1NMkn4bdYqmb18tswVbxGVLATYoRhDBmfx+IsBsS72JxADTQjccWFHZHSiCh6
Bu6qzUVxoNDGaBnahp1nb+nSa+MQTeWIbdL/MHeFvT+HT9AfOidb/7Bvo61wygnR
AyzYXtaUw7xN+epRBSGXnN39iQuxoTbLtDpU8P3/Fe7eYLGDD1dGZQVdX6daOg8U
gPhSlcFllHg5EVCs1oAVnyFL6HivF1aocFiATVW6yaWvCGSK9OU4KOV/5vl4/2OS
pUoOhYedFaXr+iSsSqc6mdvIpxYJu7cpSJ0Rc+8WrwyAISLkBFWDqr84d385ty/D
CeuwsWlhKcbgd/d/+tKF9LzqYPAP5gIVSDbW3lc+gyoTSWMXLu0/03T1UkY61Gkd
g5i2wWg94g2fgpktOF2gBNEP7hZVG/xG+dNzaSEZFJIEgV0L/0BOlxIxCq4/1mIL
WneUMjsffOBQMS1mzc+Yycsm5tDDIGk/k6zwnRWEVfSK7xKKRO3VBWpn8jXoWyb7
YEyuecCNXBC/3X6x6EB4Ivtg1CtDJjs9XmyMbGJQD+pFTPceVGOgfGLlJ6AeEM20
4LgVcxaOTwsH1f5oBMK1Fbbq5+GdYi9opQgMTdMQQnGgh2+AQTnRqz/djz+QDH9+
gCqlv4laeCa55Kmsj/Zs8SSngTBJNoUGx47vqCEY/HOOgfJ53GtYs52vYPrQVtAC
mDEcLNs3udlYlla8P0x6bm6KoCc5+UnDrfnduEv/xWZRZPDP1eEk00iGDcM7KRZq
0VT9PN+O0eKO+t9d4Y279b3A8h8WuM6NElFzYONj//E2k6hY5RTVeq0TlJTa3BA6
WchMqTJ8bZWV+hR4SV69/C6/4Qa55zfcWMynrO2hy5aa4m8u5BML3w9G7yUUC7AX
OQ/1EgOKi+aDwsVgqjoDRqn6S3/NrrCsfB6iGuiFXIkP02MsUBsrtBfUldqXC9UN
Qq1o7vHuJsamKf6qB5gDxd960Y1AJu3PV2OtdXY7wr1lzWo/G/K6K4nxhQguu8op
s/anSW9rE0wPmes2n7jBLg3JzRI5ECaHaPYFj2YpAVHhwKdEuEagGHt2nb3DNJLW
DBPaS+q0473ixWvTO4FDoKhbhxT+PLwfBz+RrQ2wgOOuJoUOKkTxfYnxMiL2oJ71
hJPUcLWjnIujFAumrAH01dPMXKjcnF4xE/6ItWsJyjGADEqMLSqutyPHoTADviMQ
JUJmbRGM8DBcyAMidnMfhmz87SToqtuN8XbB6BRY+t5w4qqNvoEvAtOfsQYbIbXi
xdo9DJlKGJEnQBgPPAtDWX52nL9vj7QCxAUeU8GFDVPrvWLQifER7+L3UuKxWbjC
fyDaPwjxm/e41di+hAG9HWbApYj5bj2pRi9QoZVKb7m38ncq70lyq62ujs+cTLjc
9eSKbhgyckY/bvYEqi/auj2a+5EBtfyiYJbKLYpnI8PxLvN6wc9V4Erowp4+d0Le
jZRjp1GwTAm828dI4cavQv4EiHGuB6kai7+H40HbC6CCV6zhB1BYjobBMM3B8g+Y
+5iQMozAvHXuVdtZG7x8MibdB7mgfjHTW9lGfVPGcgBh2kEQMOjNOkA/XQ0fqq4U
K1q4MBHW3iYYJAEIHUmMZYUoKzGmWhMUwa7FfZgVDK5JWKO49AE6P2mLO+oy92mE
OXs7H9nMNcADa4jWn/yfoas1W0aI4uwqqONb80TUp1r8kMmqnVUdJSHGmYEBS3GE
bNR0Fh0nRBrFSP35l4j+WXrbFGURCE8XykElDDgg8lZKQ4O59xz2MhOfxKrZPNH1
ahEHKbi1P1xi9GXRF/KWGPRqBK/P33YSBjbLM8AGnL2yQjXY6Qm+msFdOdOI1N/l
f6r8xWyHTo3sXAG6UgiQz3ita+qcStks7V02amCm0KC2MhIapXp5XbBTUrLuILqA
USXvWF7S8iN9wCC81y/+EPRQImZbcOC6MzeusYSI4bzmCDZIalaZSI01kKwsRfPE
8xRRVZ2XBeMNxxpIEyhx6CV0xr+ujREi6kUWdv4BIZFbYogFoq++hiRZGpYPHUfm
rJT0Sk6ouN0BPOET0Qvl418W7Ox92MtWu/f4/8980jtPBT0ZkTnLlA8VTgNwyC8x
pWZjVHz6tzhTqPBhfqECv2FLfjJ4ArjU1qJqmGIHFAofl7I8j8/BiO2IoirH/xUM
PnuRkdbpmTKVzwKpghrHrqxbEfF4J/sGKXkoXKR1cteuhHVEuduHpPGPBh/HbBL8
BqKLRz6NlL+MR4sLNoqOrvc2J6i9iPaMNDtEOl/n3DSCfnYM0M7FIdgSRxlT34ba
Tu9VK083tuNpCEYNFLC4okMBl4Q+kCL3g3LzYvY4d3rt11BjY2IbDePhpdIWhMhG
wu6pA6HfntHou2s0PtkooXBI1tt7LVMFe1wJQNh37k8wFkXyCj+3Uy2zub1X9kcb
NkgsGsqzDCFE3nHcBnutGYGkluCfmQmL1orbh+naaoD8GsKxCkbxYD89RVHHChIX
hjxyGGJIoaZVsr/nPPlFz6KXUecg+yJP1O+FalBmdEF9Wr9lHe4EeE3OJh0LHF6c
yzA9bV1e1LZ0+OEa6Ec3Ul1W7J/8tVdgjN2Bn+Fg3gGyjQrSeaxay8XoPkWao5O5
38e+hCIiNWAS0WEOmDDWzxyj8kVbMLx55H9Cleehr4iuFDQnuVPZWR99/lePasj/
wiFe7NzIUo8VFOmVbKpJ43pXcTmeRG51w/o5o577Fex5Z6GSUp7dp6snBrUDSdh4
MhBAIzzKEPNkKdBm4jLuqfh8yKj7NOp9jIRxk1kl4vf7YtaJ1VDFMrFPUYbSfnsF
CO7laYNW3zLl2Qp9eU5Ou3Qn+OabJoCvbawG02x2jxPrHkw7/rvKJ5X5E11NHjSJ
J1v24LPa2PmLPxnQkJybCVBFU4dpFux6akxktIqS96JwDV+Foc95i/2YPaO0bAur
d7qLOPw4qGGdXW4uf626HqvunUUjALd5roNI7hz9DuCbgArRi6POjKXamtFWME7J
t+2QfncKyLiLTUxx3fi8x3C8OEb9b+hJ2lA6Lw9BtSV1rPU4qFAC2+hPkZ38d9od
LBCxPZ5xz3kWICkLTJuHJLDuy8X/m9O4cP0x9vodOad38bdKNv8LzIAGJHckpz+f
57/SAmecrrmQAf765phNEasx88bko5siCvk44l0cJKa9mUlT5Y0EmCKIrU7zshZH
6vA8Vy0jAbAx/L6LI3RC7uIl/+VP5JTJj41vNc4Tj96gEWnfjTPC6wpNaR289VFf
MTIK0yDK8DPrQwQWSTwI9htBGg3xYksgPG4819kKFsznKO5q2QxVFcAzPRotQFf9
r51VqULenz1DLjVG9P4ljVRLiHQq1A2hevvwTglobBCc6cyPCx2oVkiC1b7p7iI8
hLZne/09EAQpoTLaxPbs7Gfk63RiNm+EPcAmAT0ynIAp9iNfj05K//7qN4rCe1AV
KE/0lT5rJ2lPgAmMoxTYV+jxvR//kBwYDoLFkgGe0lE1LblQQwzQDV9ME+VrhWqA
j850iKX0OcK6hB9Ct76DbHLHqpowoYEsXvcqrCGs/K9vcrk3W0s2NxZwIFQVc9Iq
ee/lPfZMw4BL/LHH62nDp7qv5ITX+HtxaxLOdQ9BIQ7AyzPic+YQ7vjouYXlSro/
8Y7alqabjqmR9GNsw3DrZkZtv45+fX7MoYpPlrnWTn3BrWuGFfrYboAO1JsaKt5M
N40jG7UmGh/rWthcRJYklrywWPq/paHt5Zb6VBQj+MqkWzDuQkUlsR2rTEN/mQ5f
RBSOHXxL1pKm3UDhzj+jLOONyDuMVFXRotFufpNE2yLkZN6zPjSyzPr1SxZKIYxz
ZtkSe8gtze52h1U4i3szLxI+dtguK2t3nnh2l4J6fIcA0IVRIjIGtuaEbv6keyqv
2rDu7qwQMXnhWk4qW9bUuPNe3cftoMozcQ/xw00zXp6rHn6RR1EYvVzBTNGlPYKi
uPGg96KGpcuDoSYhQjKy01n6u9A+waBQ+TmfIW1VVmXssgSvmuqxx8YAeq0vti8s
8bEZx8ZQ/tXLNjU2ghP1ZA2or9qvY2laFk7q1Md8WSYq3meLD0u9GoyXZ4jXM30g
3ZGz7T64iyVKfrTE61Nd5hOrPYr6ttMxR4P51rldFqRO9ZSQ9bIcreZ1SXnEaysX
eE5DQTQeHeMpXPJSYJqB+CpYtDD4vyU9n74nFH4O0lqM1CvVqyII68eK8XsUZh/K
JJCcipjt0gRSA6rQbLzIlsqdaXWj05jSgc2Ct0t8kteRklIjhzLNV9DhLmePTeyC
4Pkr9JozGg6a0sFwofIiFkAC5zVVgrYqhbezz69eVyJND8XCx2aBswUJA7tZ1Sk6
u4lY1ng7+ofxCumihV3NEUz6bDXGbyaRD3IfqTqJqH8PYrp+1GkkJJ1v/GM+D9Fm
ddlAJBzwAl9e3vOZsSpIP3Dtlcei+xcfJk6Ze7gSF4PTdkeFREjy66/7t5hMwEY9
wBEKsxY2KvC2QRLRKi10bt2FRf4mm887s3fqoaZKKoiANYAYcV3uAeSinP/Lk5/f
bmFWCJnQGRBCEvnfbtACpaKODN5AUaIdYjjyLQPyY3jDMTPC93J1sk6xYEr7Azlc
lJq2THY7HpPF8NjRf5j6FbyI4pLNDDeaKrbTYQsC0kH8ds44qkrkfvvQmNhBpLXt
t87PWlt+3Q1GiHDHTGiF+P3X9iPhlrFmqMMaKECOWVsJFblIQcIxsfqtZnYbUG4W
dq5IooxIeuCdRUJRjd2JdnEhQuU+ediSH9S2HBQ6JhKQ0a0+XdFw287O2wlDzXCc
Quy8t+3ZD0Q+qUnoGj+xxpoIiHc86Fi3HAV3Bnm82Dxb+WOrxbxt2vvRTOyeYJWA
v43y+V1heriH/Glxc9g/2QxjDeUb9Vu45nuSm9+EISHyPC6F9L7atGZ9AOjYcNS8
eNkHqOBCxIVV4Y1K/KFjZLCoGGR718Y9S3X3GGc3aTu5aOl/mObAFS+lVyd0+CjE
+d983Osz/V6VRllACWDpQa6bSpssEhyu5EAzvkCcrnyoOSURy+V67YtFt//tctVq
+X22OS9pK5VrffmIKFB/4UDsXfsf4hCg2E5Z/4U3d0/n7XCA8CqoBB6zUls2c6BQ
sTaVH6fODevh8ca0iyCvgjIXKq9YaoQpgkeNKslg12q6P7yBtCyONzYtgnlHOu0i
bWxxxhNUF6+K79/Tr9c2MMl/ipHrSEeUl9VsJj+JSLxbftOx82ObNPi7rNLWtB/8
YDzq8X0avHgjXWjg/9Yz4sG8pr1Wf7FfL79nan+l1hlhgsUPEeIp4D2J80Jp/KaV
vgeEZ8Wd8cA8CS79QOB0P9qf0QQ/6eeZOhImSkAcyrNv1mgm4mWrpZgujw+WEwv6
AGdZdJvK2bgrzgFfKgNV4uXreiaQ0lY9hU3cdpyJZrdpLZzuuI7z3bEVA7DTcCbA
eyDJAZtVB18lmr9UVxrysN7ENVbX2LRIBo7PyidHk0xkQnIAgAnrkCwX102jpeLe
YNDxzFaz84unGuCBqwQ/eoLTZQdHZAQl40UuSR/dCiIDoq0TSXCmORR9VO4xYaps
+RMZ35GiW19svny8jBMKm7NsRi31UuLsjOaIcBc3n8A5tlSHrrcAzmy4spZw/PVT
F0N4UwSQxuPicjPzJSKEDqLcKqqtmXwDcX2RgaMQSgPsVPDrivfXgPfBWVGsVd+5
zd6g//rZVeNhlEJIT3ZnkYoWAY9ouDrhdDs+NePR323UaXlJeQhkByuZd4XAxoSS
Qy9n1CDKA0Cz62h8ibaiIMC4Ynz4ENyQKRBbyyZzyJ0Pe3hlcpGAOYAVW+lDtCe5
M71D4WFy4oXkcXNloZZf0nGBgppRJqaBeac0UKAI+GGcIXiLMYs0CW8KQSpaIKmX
mioUQgibuXE4A2MaQFN5+A66rf9wGyFM6vHN1QNVwrz9eyYuGd2Y+L3sbgczy1v/
0z986cKy+3g2dsldCMQTLkVM+REHlO80+Q4z+puKUJuOSPlGPmclpgx7MD57R6tZ
JefYOnWUkDMYp+i1q/11crcUPw0NkFnGCZOJCpMMrD44eM4hKlc9OZdctaWMMmte
HP+jzT7DaIBEoqU2PrLFoMWu0OG9ZoRGStsQFf9MwioFrQhyAD2A0yr7jk3qDAjQ
mYAZlJhAeTeItfBLT4/RyWvzZtjPgVwXokl9pEIILXIzQBwdywH8QRRiD/cAZQ7+
i7CB6rSy5IVUqaNLNJqG+GMMHBkROa2b2MN4tY40qKDz6h/A7t8X738VfPW/dlBy
ztbvCmMIL+WrvHK/r7i2/Cldd1TjZz+seDnUlbSL5KpCse1i/j2FV4HbHV6wfa/6
8E9iqCJm3lnqN4u2p5uTZ6Amfj4NTjGFeRTh9JURnRNFy0bJB9tOS3Vt1RoMxu7V
oSMQUhDhstAwUELmmntvvxVsdrc9sORdT8+4YfqVkjbM+awXiPf+O2f7vuvIdtUz
jlhdxMkzypkB0w8gemxwncPI4zGnzvDT5Vm4b02r7uIitWCtNOIdrnUPxhOzZoKL
SYabobtWsBS6MMX67L6DI0+0L/LzWn9mZ48w3arKzBALAVUwlUgbX5/uSMgM+WJz
pyzcxO7LhSp3cdnpODWYAzV/pBBoWUlapcCb+3DphorNHPxiXdsHqtbKT9wlMw4R
wpgRiKCWkTo8R3UadAtNjr1q4VVShtjGVa/dWLEnKEoOYt1xI8hmVQYZFZ0HsDM6
bSONBbAEIIo3/hPkOlK8iccOgQTZhKLANPcwIKC2fThBlHG1YYY7wrN/cVBNsDZO
ZsdC2ezBpbHFVF+cCdnp7QFfRtflqy8V4wP0WoLHNVyYTX1hIQXRQ5mumA/pWY4H
gi1ZKCqbHtpTmXJkDM8V9j4AZ1DpYNXNjpX7ufY/guncBW9aZ9joK+6hZ/IhvIxP
5Zhb17O9+/zyO+o50SJOIl5KgDEVN5bW8zLkeHQy58j6R2AG8Vzv1FV1uG5EXrfI
I8Xk9RDRxObX2SB7gOqltolT2+nr3W9xOG3C078FYJ/QQ2KPQzmuyx026HVg0p+f
ParXSOxOTXhH1JhlWZSPh0KaTyzDkkKJk/Y3QWLRbnCdSZJb+rpUMt8IZZc2vnXh
oQ4obuimzLJ1vTsduaMhpP5noKFTw4f+/FcHndQkOXhBZ9ochg8r4gmvpc2GCazj
oFGSnpKlUocqypopTaNF8uwf1xpa3hMZYSMZ0EVlVrpCzpLGFlNIrSx21wbPL/FJ
Cp0VuA74PX9sv/JpfGc4AOnEQQytG7y5nTeh1n9xj5/twNKMuVuBtfOQvPuyPUK0
zFYt2qOB8uYWlH3gT4iPAqhh7Puz7TaZPstbOczj0d3zRUhxArMdLqTn48aF8/1m
pYLRfJRkyaKxkwyMvSyrP0eLYK3p1r/vprWr12Q4relIxWhqPEpxShqlblcIcxyQ
pkZ2iff1vXzbJhC5ONiJ6/TyouUd668DzJyt8lcg7WPeQ2jks+Fq2vrPEMAjs+AM
yIYm7ag3K5mH12s41shVnB+680rvEobN2At+3qWA0WdPdd1ngmYCTQQr33d+UaEn
V/8Zerr+NGYw003+zHsapMAVOtwmzij6d+NHZ++FzXRyuHjneS2dvSmdvLqeGm2d
OrhGM4mMfli4mN1+MDDv3xE6Hdf0Y89EeM7+rZLhQQhep5MC83Rr67if1EMbWhL9
N8B1lqdiUOrGzOs+fSf7oapBufBr/khkyT3nriiIpbG7VTi0DPtEZAWsUTw/NQT2
h/EVQGg3ZNrQHJSOZ7VOydiTG4lodG3puz5VKook8IQ0c82OY79HyeFPH5YSzL4m
PQcLziBlyAcne8i8qCLEEPwxsdekJtFm97TxmBtrW6tx+lCohBN8mhfLk3cPicQn
MVBso3MyOcxuE1xL7FOf/w+h+G7vuW5/fHrEwzaobua2yK5FbZcOnM3PDihtWXUc
SLhs2AdSJgol+kajh9bHopspDvUUO4q2LyfBqFTRFwfi7Wn6gCk9/RKvW5dMoGWA
tRPwV8RxXuaTGENXyaIvmSthMXNaMZT4LFlbc40WV/ZidAYp+0FUPqeWAOwrqrJ4
TF7jzXi6febk4E+o2Kf8G2RRK5og1EEgcqSCDodhsLbr89Wjts+/GFwrZEI8CntZ
Jwi0YFSnQTW+SiOn+stGIVBMtOMqkztkfZQA9Wtp9b1iPMrhJYwZPo00NB5AyITB
irVc4MJbF5dxVvll+umxHLdRAvMOgs6FoxhdPKWVY9OeG9JDiqaxM89cxbi9Ym9P
L+XZ5mH0gb1257JdxR8slOs3RJmEs/ed+MQI5ef4CZjt9JuMDaRuI2QcmTFhPsaK
WZQwsDdpyp4NmzSQn+/Sn0Bq8QnYLyOGHwzdTKJN3T+hpP/4qphmM0i/4UT589no
unFi28ApKSil5AZ5eFNQIDlhEYTvXx4+yBlQ+18Pie89z8kdutcuqYzyp2vDxqDi
jbOkZPjSgJkeyqD07ANt9zJ5fDozrHNWkxKayCvZyLHhZwUKpGAejFQy73pNKzcD
+hHlAU/GP0W75DvahIIaQwb6eWdDvDcXfJ2tWuOcedPpwJp10JNp21vRU8FR+97J
ywP/yPJz36zrsQg04prRObL7k8o7ZxOQyUVysyBlDKAagvTqVeuzU0flgqx0LrJq
rf7WzoziFvMRtrX2CmBhush2Wy4nyuJofMdfZ9vl1yEjbd05I1HKP4/FIk+9FMa+
1CCIucPuDx4/tM9m+/AHddlehUZtXkWYAbI+FtbX1V/xmHzzCd7nAGxGHHAfU2xm
/ELXJOttc9O7UQqDG6+HObn6GV8HpqjnnW6Zlh4OOvixoRCc2KxAlQ4UiUy1LiTW
Tooi4WfOom9Uv5BMO4HFwSgfMeaP0QsHidHq/0amUinEW943xAcdVlotyh0n4ppG
UcEaIAjRkyKOnVqa4iAyIuK0F1MbAeeMzDXYP6/TmRiugKjG63Obq9aVmzkvB8KU
jg8hudNRfQYi1ekmXS6GjaQB1ZGtGj8MCBMw8mYgzEr5Dw8WvGTH+N+Ctq7nrQEB
8M8+wY99PS9bZQEh5f1UttkcZEVhCQu1ubnyRLVHu7YTFxnws1fAbmAeLYpFHc0F
apmrG+PgmMLRp+RRLlpBf/lVCQodp/iawVvgF2LXWsX7gSmk7L/jcxFQPgGdXi5i
KKC5666C2WylyrvDiIT5+Yz1RdVh6nmnZTRuc9S054oLvI7SsWsCbEnDsITHY5+r
1e7W0ciQPruwntbnOZ2CE8X0rsGC/TcHOD/tUhgoXikDXy/3BIPr7DpLeLX9a3fp
QPglGcn4JSLFDYHV7qwfYxiHxPtieY5JrbFfqDge4NdFqOvpm5ZbF4lYvPywcYfa
mPc5u45j84cFoWTJkTlL2lDWEeqGxGDVqFUJB3FyLgh+bXUVp7zPJsJqGDawqut1
4bdt0nAgtjeLSy5VsyBzE/A/J72GuxD7883wmxgAYwObs5icxDqxM2aYxIu0UKPm
7MeFwgZ8MmcC5QLn8Mnvc1JAqzqlyqZ6EoSlUnNLau9SOHZHDC1AvkugahiKAwmQ
Z/dFBGifnFVmLXs4NLR8iD+DkGES6TIx809waXKGBNINjP2C834pJrI7z+5DykLS
DWqVwoQmu+JagZaJI3Wn5m9qXz6pBF7ZoIfuhJLfuy7hKOWnFe9ercpwTfGtl6Xj
PJeWqrKevmgyn9vEMyd9IsVxkTCTZu4QHIDCFfplxM9xSWidflIf66I3N9N4dxsP
+nuORtTfEwdwuXnywyltgG2owymVvxpS1BDkmFo9zInSfMBhND3v2BXQ81JxDOi5
2bx75028zllanorRp2mDiUR81g891undPnj3QdiDyvE5HIc/rl2IdxUU7rM2DrUj
Q/SMbbtM0aB/qjR7Dd+0wg==
`protect END_PROTECTED
