-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.0 Build 156 04/24/2013 SJ Full Version"
-- CREATED		"Wed Dec 04 21:34:39 2013"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY system IS 
	PORT
	(
		inclk0 :  IN  STD_LOGIC;
		UDCLK :  OUT  STD_LOGIC;
		FSKDATA_BPSK_HOLD :  OUT  STD_LOGIC;
		c0 :  OUT  STD_LOGIC;
		locked :  OUT  STD_LOGIC;
		RESET :  OUT  STD_LOGIC;
		WRITE :  OUT  STD_LOGIC;
		CONFIGERR :  OUT  STD_LOGIC;
		SHK :  OUT  STD_LOGIC;
		AOUT :  OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
		DOUT :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END system;

ARCHITECTURE bdf_type OF system IS 

COMPONENT dds_config
GENERIC (FINAL : STD_LOGIC_VECTOR(6 DOWNTO 0);
			PTW2SET : STD_LOGIC_VECTOR(5 DOWNTO 0)
			);
	PORT(CEN : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 TRAIANGLE : IN STD_LOGIC;
		 PLLEN : IN STD_LOGIC;
		 PLLRANGE : IN STD_LOGIC;
		 CLKMUILT : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 DFW : IN STD_LOGIC_VECTOR(47 DOWNTO 0);
		 F1H : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 F1L : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 F2H : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 F2L : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MODE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 PTW1 : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 PTW2 : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 RAMPRATE : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
		 READY : OUT STD_LOGIC;
		 RESET : OUT STD_LOGIC;
		 WRITE : OUT STD_LOGIC;
		 CONFIGERR : OUT STD_LOGIC;
		 AOUT : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT dds_update_cycle
	PORT(CLK : IN STD_LOGIC;
		 FSKDATA_BPSK : IN STD_LOGIC;
		 UEN : IN STD_LOGIC;
		 CYCLE : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FSKDATA_BPSK_HOLD_CLK_CYCLE : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MODE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 UD_DELAY_CLK_CYCLE : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 UDCLK : OUT STD_LOGIC;
		 FSKDATA_BPSK_HOLD : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT clockdivision
GENERIC (division : STD_LOGIC_VECTOR(5 DOWNTO 0)
			);
	PORT(clk : IN STD_LOGIC;
		 cout : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT pll
	PORT(inclk0 : IN STD_LOGIC;
		 c0 : OUT STD_LOGIC;
		 c1 : OUT STD_LOGIC;
		 locked : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT testcore
	PORT(CLKIN : IN STD_LOGIC;
		 SHK : OUT STD_LOGIC;
		 CEN : OUT STD_LOGIC;
		 TRAIANGLE : OUT STD_LOGIC;
		 PLLEN : OUT STD_LOGIC;
		 PLLRANGE : OUT STD_LOGIC;
		 FSKDATA_BPSK : OUT STD_LOGIC;
		 CLKMUILT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 CYCLE : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DFW : OUT STD_LOGIC_VECTOR(47 DOWNTO 0);
		 F1H : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 F1L : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 F2H : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 F2L : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FSKDATA_BPSK_HOLD_CLK_CYCLE : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MODE : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 PTW1 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
		 PTW2 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
		 RAMPRATE : OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
		 UD_DELAY_CLK_CYCLE : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(47 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC_VECTOR(19 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;


BEGIN 
c0 <= SYNTHESIZED_WIRE_23;



b2v_inst : dds_config
GENERIC MAP(FINAL => "1011000",
			PTW2SET => "111101"
			)
PORT MAP(CEN => SYNTHESIZED_WIRE_0,
		 CLK => SYNTHESIZED_WIRE_24,
		 TRAIANGLE => SYNTHESIZED_WIRE_2,
		 PLLEN => SYNTHESIZED_WIRE_3,
		 PLLRANGE => SYNTHESIZED_WIRE_4,
		 CLKMUILT => SYNTHESIZED_WIRE_5,
		 DFW => SYNTHESIZED_WIRE_6,
		 F1H => SYNTHESIZED_WIRE_7,
		 F1L => SYNTHESIZED_WIRE_8,
		 F2H => SYNTHESIZED_WIRE_9,
		 F2L => SYNTHESIZED_WIRE_10,
		 MODE => SYNTHESIZED_WIRE_25,
		 PTW1 => SYNTHESIZED_WIRE_12,
		 PTW2 => SYNTHESIZED_WIRE_13,
		 RAMPRATE => SYNTHESIZED_WIRE_14,
		 READY => SYNTHESIZED_WIRE_17,
		 RESET => RESET,
		 WRITE => WRITE,
		 CONFIGERR => CONFIGERR,
		 AOUT => AOUT,
		 DOUT => DOUT);


b2v_inst1 : dds_update_cycle
PORT MAP(CLK => SYNTHESIZED_WIRE_24,
		 FSKDATA_BPSK => SYNTHESIZED_WIRE_16,
		 UEN => SYNTHESIZED_WIRE_17,
		 CYCLE => SYNTHESIZED_WIRE_18,
		 FSKDATA_BPSK_HOLD_CLK_CYCLE => SYNTHESIZED_WIRE_19,
		 MODE => SYNTHESIZED_WIRE_25,
		 UD_DELAY_CLK_CYCLE => SYNTHESIZED_WIRE_21,
		 UDCLK => UDCLK,
		 FSKDATA_BPSK_HOLD => FSKDATA_BPSK_HOLD);


b2v_inst2 : clockdivision
GENERIC MAP(division => "000010"
			)
PORT MAP(clk => SYNTHESIZED_WIRE_22,
		 cout => SYNTHESIZED_WIRE_24);


b2v_inst3 : pll
PORT MAP(inclk0 => inclk0,
		 c0 => SYNTHESIZED_WIRE_23,
		 c1 => SYNTHESIZED_WIRE_22,
		 locked => locked);


b2v_inst4 : testcore
PORT MAP(CLKIN => SYNTHESIZED_WIRE_23,
		 SHK => SHK,
		 CEN => SYNTHESIZED_WIRE_0,
		 TRAIANGLE => SYNTHESIZED_WIRE_2,
		 PLLEN => SYNTHESIZED_WIRE_3,
		 PLLRANGE => SYNTHESIZED_WIRE_4,
		 FSKDATA_BPSK => SYNTHESIZED_WIRE_16,
		 CLKMUILT => SYNTHESIZED_WIRE_5,
		 CYCLE => SYNTHESIZED_WIRE_18,
		 DFW => SYNTHESIZED_WIRE_6,
		 F1H => SYNTHESIZED_WIRE_7,
		 F1L => SYNTHESIZED_WIRE_8,
		 F2H => SYNTHESIZED_WIRE_9,
		 F2L => SYNTHESIZED_WIRE_10,
		 FSKDATA_BPSK_HOLD_CLK_CYCLE => SYNTHESIZED_WIRE_19,
		 MODE => SYNTHESIZED_WIRE_25,
		 PTW1 => SYNTHESIZED_WIRE_12,
		 PTW2 => SYNTHESIZED_WIRE_13,
		 RAMPRATE => SYNTHESIZED_WIRE_14,
		 UD_DELAY_CLK_CYCLE => SYNTHESIZED_WIRE_21);


END bdf_type;