`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9CssApn64BjXz1XhoiUUzjfluiyLF6tsnN/DKkteTfiWeGn3nErFXmPY4Wpww05k
zXbxb3oyB1iS84CVUB7CvA5JLaa5JOyna1PlGoDjO1f6zxwSpfzaM/1nfVn1GDDH
5Yy+GufWc771H4ST4lPb9iImc+UPJgyeOxzZYeGhc3w5T8mcjlKRS8E4O2y+PyJU
kzcf/0QIf0MqyyrsYLi5RETEdZ0AhSSO7XKVyQAl0nxqgtnjHu4uuf+592geOup1
9mPO2lxYswwh+JnNJ9kMQrcfGUyf+tkHywZmhh0IzDOdh8cYENk1t5G0aEGWuK7b
2lnaUEjIiXg9JG5vwBvNM21KxAZWFvNhliOEOeNI7XWo78iuuid0lA97OTPg6dAq
qdnzlEWNbAKrl8wdbpniy8epfrsqDHc5EcaIUiPUatMJdHm88O2YwNmg0nVeeU+M
C3h9baVCKsWelh1AIDacf3YQgR/dsDi8hCco96GPHDh3zlUg79vNfo2ddkLzF72I
fu8IaMisj25L4Ksypo6ssi+RHzEqhRq+JW9abiawG05TCMk5xKRPzshoCioXzSrJ
y9TpI6WDItuh+xWn2s8X3PwCI1W9LGQx78Tpc9EXZGC+MX/Czju3gX8SDM3RidGr
5/CqgZb8K/ou+RV+V1uZF301eL8B46gXPLuMyHgbgctWh4FFly9skv5NgVRyEiMv
wz94sazeKurVhbacgsygEr8L1DTlCLXqs9fgjV7yWbEXR2FZdKj/ZLGqcL8bewBm
hqIYqLAJZRI5Qc6dXvkxtQUIfQz43bhYimLd2iC/s4Y6LzclBCDn6hmSCHIvoEoU
4bnzzrB0O0yKdQRfbPaMa/dKYZMAy/OTx9WYFKckXe81qbrwauEs2XErG1V+xV4H
1P8VKhU+CT7D2lSn9ZCnxdbG4mlZY3n4CWQw6WTccUYhUAfUmu7C2qhBONF3aSyk
hitVmI78xKtU8pLwN4l2vIWl/HIe5eZLdtj+LnQHTixYY9aNi4v+13WAzJY3fClJ
OISrcXWzRBY7FMdWiVurEAtyDVP4fpNNflrVKRpncc2Ja6zXclPj5xXEZjAvKrk5
cP/DgG67cPJiZQDgTJwznHD+Q7SKDJuU8FoMAXworncXds/UaH/szFzlZfPf5LB+
66cNC9ljVQyf41AxP5FodBS6p96z7Juz/YMVbviQ12xG6AcXOgFLZOS1WiTQroKN
mF/YE52Mkozf7st5yZ4ps8L4K4O8MHdZ/QWG1zVb8qSPS2HVMb9NnT2WVToEEAZa
ABYe3A77AAoSkpC9eZoRx7QxIbYJpXKMczRJeUijOKq9hBYFmQiQqZrWG8+xA7Th
rjVHZGAM+AlTEjjF4KOFJjJ3RHzBaCMiQ+HeHgo94eepg/0LrOgvwCBLWT7r38Dr
9Ek6SkE1DcNeCkvCzpFBKmimkE/uZL6gqeeSI6IFefnVvFL6AbCYBFB1Kk/5XdQ1
JHpeos2ScGiNvahhvR95Wr7aJDBwkmuf/B+60mSB4031EVjhleBT3NCJTIfijr/4
d7aTwF5tjwyKhciMC11kTXNEhUY5z2wKPPU5i23f4c5KlJ5jMh7sA8b68ZtQw+wx
7qAqvieMwKzMGKTn/IlwvyllG0oNcBaWidQqR44c2WRrOK6XkJjuUpfQHRN4idyB
/jlcMNDgyp2IytbrhtWG2HR3dTD6iY3eJ9WOMaG/w8T3sonbWAwX6J/Q5wHRSbUz
ISeTzZInDQ7djvSEz9e+tIZx+aJX26EQczEDAfW7l7pu2GFDqSSWr3Q5gGjH60ll
UsPM2jQUiwowD92jli5iDmMOfVxIV2PN/IlgG8U+y4gkwsIjFD0g/epTY9SWjdi2
BQK6zZNVlby0Xpck05KdMDdTLHYhX1763xlKObw73DgvZ5gB1YZdtDcLIeM9CfhX
ZbRxo6HxXLCP+Ghp2xrMXCJcgvR3l+eCVjTQTJbR6WZLZGJv5l0SZFzInGjNhZR7
FdsVMn66g5ivKC6gbCqWSHSKNfr65SfExPDz87UvYr4DYpJmZECNXxSr8x/+X22z
BP9FDR+YnuaPvHhaIa0UM3ymuoA+uGqMfyzLR3mwwFOjgxGyA88toowsOGWRUnS5
okC5/UMwGluU2L2CFss6d1i70jO20kpJTZuT/TXLxh2cP+sdMI1+t5c0Ot3IPXJc
vHRnu2STZxBb4Vf8wSJN2xCUr3NJecsqDjrTSKKplUe6jZSssanO80xFRW00RzS7
1DJpxg2tD0Ze3kC3ZOFjGeBy0IOtwczi027eH0SlPr9UYPo9fnCudZVw9yjot5lT
oQRg9vWBP7Zk4+bvqA+Rvrbuq0HG9XgHBf5jqPnDXUeggGoy11BJWkaku7f7XIrg
Nqh6Z1fql1czmaeMbEPDyEHSLgwzp0y6YSEDDEus8r0tYrsU2hBfZcsXW0zNb0u9
jSqEWJEzPlWsCEF5njcOdLVtFL9j5zBevJPJJ4l6iMLQhjxowYW2Ev7Z7z51jupX
ouMiVWLtertK4LQS0op+dL5JBwVpRMJc+r42AMD/RppX9+BXCmVjqRTFIdUJpfib
v1/K+SS+8/t/AX9OVIHXze+CxY+z3WQa3qxWHZnWLRWoAs2beWlfsd1dKA2TEL3J
1qZOS7k3rlmvg+kuyp2bAcBc65PSrQz7Wwgpq2X+ueYLWx2RxiGHQkU3lobiIs3s
xuhZhDblwP+//o7tC6lpZq2oRhNdzIN2SRn89aVV6qSx3q28i0BwxWrnuYRdOhQ6
zdGB+SRO8TFjkk6lXZmCcI9dSxnKBjbGQanWsI0kwG5QEGaPolZZRCbAu8xUI/TG
WJjZM8Al/OFIe9FAckQs1A1eovDssYex/VsIfv2FpL1Ozjk1t6g5pZUKw20DgjPV
KZAGBALAGBgL/TZh+2FyLqE4mNUFlmVuSgUYXuaKaKsr9bteuudyoFX5VVcLhb8Q
LtmxouArsdgE5FdBvknX0Y0PPBqshU5y/0lqR9JoZGCjEMjeJ8tFtY8WQs+h1jY9
NhI9G+TD/PpIuF/HfzeqQqFZJ9RZe0Qt3t4VYZMpenFgod6D6YqWACwFR36F4t7Z
sF8+jdkNBonUqyZHy2IEr4s3iWl4AGuyvPr0RgoOuHjLAltaS/cLQ3n6rl7AbmNx
Y8upLw0fEOtI8utXL8lWHj2os1SVfP5/J5vZkEaXhpU1KS3jHAXRuve5eYfn1rBm
N9XUTbwsN5BgAXtVKtEA/ONlkfnMRozB7WvhBZVRbYUqpEdrp0oTe29RD52jBZdi
Z45R2fMW0OilpiTrdloV+a8C8CdwH4T13bWZlwoAkGeVPOexUXlHJjTo8gK+bIuF
d3F435kTlbxiScjKMSikVkqOcRDVq0xTBY3+hQ85JofQCEi6WxggA88zmAVHQSrZ
s2sn4GADRfVheCtlLQtzMgR6kIRFhwJktRxLl/pGzn0=
`protect END_PROTECTED
