`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k3eiHEf2JwcM6TUMnDSvAaD6WBdGlyCSw/wm7gUFroRivHHNpgfpYT3APxRWSptI
MDyb8IWceRENovtYMJeC4walaI5/p/v9jflZV/B9WVcsxLX8fDLefNvO9FuWlDla
P3OWiuWvw9lo0o1FCfQTxKgYV+xxvAWX4eT/s2J32SAwITaPt1PSttP9a6IxSLVR
28/AVJgvSSZvB+5runi9Co+t4sgpbpHi++om5M8FnFNi3+TyLmTCwZNJMtU4Nexo
BynYkEGq82UsFYeUXI/SdcT4PlWHEONJ3KFVJ7OCpdcNYYoU8uYrvVwJ2Msmhdnh
/Ifj200DHEnTIkD0NeJWVkjEp9m31AsDbp3w3swzP5cFT1teMN4jsKY1NezrYOc0
0u00HCI5iokILEb92DY+4LQADCyLLO377kOYY95QLu9jAXvJ+4sqpcW5m+hKzAEq
BDXxoTq6HXpsFE94xPKkF1tG+3jrBrCBZgMAat132sbcky6KUcTxgBb1LFz6NxUp
BW9UKJzRp9M6kWIQ/pckARdxkNt3vvmMR93ZWZLNaqb3EafaOl2gcIHnIprIAMKs
+hoGYVlCcFF90LEGb634x47gq7Qmm9+sJvC3+MqdG1nZPc4MPFLS62rPZCIN6Vco
8JNqnkw3fy6Ie6lEjsKToBs03hsJMHPcyeVE80oYaoQKbw27bwLe/2R3qPLgNDJP
qbsQ/LZdlXBa+Y8JR27COtVfvVDlJzwmOnQDEKdX39M=
`protect END_PROTECTED
