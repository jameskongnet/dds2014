`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rzbMvIHvAr6oqs8caKO0f02voddN2qU8XW492hGQ5BkF+8QNFE/FPEgr0stxXI+s
yf/ty7EqMy+qq+DPuQBwr90VOgj3haa/IDq3J6deJHtADU3J0O7vVBvQNBBWMbjJ
eVfjGtIKUaekk9P6vYkbPLQCZWyNAsyT7DF6nalrnUkZ0oyBvUyDzu9lU1foVbJF
fH6yx4SqG0jyHQ27qSF7dpahy80d16nIdpxMMmupS7uHcozJvqehc8nth5+DWPNd
qBOKxcKFkB/mBxRsg9P2zEigr0f6CSu1+zu+Fh6hAGzMSS53h7SFd1lTEJ0SfKdW
wM4McIlG0CSF3YLS+C8gLkYrFgXKmfYy2vnh83oXVEBRlIpMObKwSqsY56I5HSt+
nBXWOCjuHw0X/Oq2ep+sVOfRSmKf4H8XVhu8JYpg+8yKe0ff84iEP6T6i1RReAwA
Cv5bpBWxxr7RNN4SvNyiDuEuOB3hwhqRUSPXG0WjXUbfXg4idjkpajcW8Ms79XJR
EcmDXvSKHLZwJ5Gf60OiYYGzxns4sTDA3QTHNYu2eqV2X30i26xKOV9jOhVe9xaf
fUGKXFhgP8lRhlEIwaKAu+eqtH962SvRHQCVlDBCY/Aditb+9o09+r5S2Qx2byIN
5kmUZjAHeR6jNBCJVdDSfRqKcX9ZgYlzjMN/nIIXtMmVEBLU9KoGh8Fn8mDaEc1x
l9JuOmGi1AtR+yvx8LCJ3gsQKV0ONViKHxjs8pE/8JwDOvX384+0uTwIWiRjZqMo
dESjbegRIzxdNVGvNgF5ZpeQOtmWkfZii/JIRQwtXaQJ9lRkb1Ftcz60Z4UimozC
XIsn1DCE8VW5beSwI3qOv8IvjHzRy3Fl8lbfz3vjdTr25I0z51SwzOuiFVCW129I
fdXe9Ik2av1uZ+ng3bSZ5P6SyHo7YgFT7bhu4iPwep/ffjpQw1RrNcPGKTxgEDg5
3REbUl2Oaed8GQ85Ignr+1ar9vGAMeyUc7ZRdp0I0jAKNLb8BR7d1M/6JBIQ7DIm
y/4PUAf+8jJBkQqg1OAlVSE/H/BKR/7qe5YtUQMBewpE8G1JI8Y+K4MMMF2Mjk52
DFRyAPSVPAnFUVrtk7LOr7qEwDjFm120L9hD0vqexJQW+rj6F1I9LkmC9RuRhvDi
WFl+KLgs4g3AfPKryNCqGZpiMdcYvMaxhdtDRqC8zhOjkSXNxrNdMCR7w1wuJ8CM
u9pbROXUF0BYwxxazBQ9rKQi8eqWfL5byn3vH09iu5COqPBg5fsBnjYRZb2VJCa9
/q268QgVlsZkoffbR8hfCICcHdVHlBIE8KLSA/cqNcRaKgAqKjmu33yIAdP7triD
AorrounDWeCxMHqiKkWO4dpQQ7B4ur0rXQqujo1lnQ9PkC5d62JehfF4duAa/fAk
hMZAJO1XI9gwIDnfa+zvlEGMa3xyPH85Qpy+dMXdzxOJGy+7Q1gE5Tzm025zLLmJ
9lyvLVlVJ67JvggoB+O5zvjGMY4V8LNfQgufJJg07nedw/vy/a6BgCjIBCr+5L05
1wKtbpXxgCd0JIkoaTDPhWB4zuVZPC4MFkIfKf5NFJk=
`protect END_PROTECTED
