`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zrxafM4Dnu3GkyYjWYIIeebw4y1Cv7ZeORB8MVqI0xIQyh8UOiO7aWI8k3+uY3Gp
rZ+W1obeLMIyPL740Ks2CpZkviGEkUnzXJTh+a8P8tkWLSig8mhlEYhfIM36xZIN
ezXJYhAbdbPcwGrHy6vhyn0rBgO8E/4GkY5NjQ3bhA7LZ/KqAKOd6cUyN7WYceBV
mmdk9GeaTKgaCe8S5DAO2Aliv6iCOyeJF3wWkwx++ATvomG7+kLzNZxqZ+sO/S5q
wvuyndkAV87Ovm7z0sQw6t2LWIvpLUpWFASIK76GryXJtgJzHclyI5z+a94i6oJR
gqU2CLcbeSUiAGENqgrgDhuJ3FeUiAnNikj0ONEZiIg3ikZoMoMMgc8fj2SphS+p
7cu3aDmfa+zfZDbFmzfcRI28YvXA9eMylJuHotOIa4kUbvmAfP88s5BSZR4eakcx
7vwFmOkG7osVbQHa3H0b5DecW8N/jFTrZEDnGevAGZpPe1ETz+An+FpuCVUnSCUw
M/2mKYxalqQyJtVCRjOQXu+/2OnPutiPnTxu9q/fBlylvnuN+EZaxX4rYfxmY/jS
Enq4vAJhAfrq/0g1FgOONwvgx4MGju5bQsLForayDeH95Ecjj94TFKSrDmG/ERbK
ZhQhdtcVjRIgKHYJjX8vIi3og2QQQZyA7e3lrdlVO+QleOY72ZJOF8uLODJ8E7Gl
0NWlo3ctcnM9LbC2A/y/h6q5lwjKwOQS52xcFD1Pl47lHcneW3G83WUHN2pKcmJs
/zVer1CgUTzAXOmS3fEO8ogjOH2zuJuGF1iX3UDkDt9q340Ql9Hs0lo68chszx8F
f1iVqoUCeJXsqDjG2mvneYOQff284QBTq5Df8gYbC3HmFLxh6EO3KLog+QpCAY9O
7vrvFCwurt25+zNM3I0kKNlIM7O/dfnwXjalpkizopDRc5WdBOyMBi4ZtUvtU5GB
mIwJvxMz5xXd/1bRoEbSi+PVAPj8KGoWcMdJ/OvtwRRWN74MxSegnem5WdGEmVrn
zx3EeR0zGA85IsnTX/NQD2PHXjT7YCWQ0KUJpzZiOUxiQbC6eWh5xliIKmWQeze/
mZzzc5jHE+jtSQtQrRk4Xq7T07vmS0Fe3V1eZbPdxG/EGJoCf3MU7HS5BtE85OjH
QvlnXGbStIm/pBM+F8rhGANbgi3eJWPz53AV7k6Jt3bcQMPMxhU1ey/JDO6ZfpJe
jQBKfON7k8yz4v+m2rDjKLVos1vUkGMdNNhCbQUlnzc=
`protect END_PROTECTED
