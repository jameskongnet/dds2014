`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hDe0/tu4jzMXubGrCBVXftKb01A/3cca6HsqAv3CN74wS2yNJNQhyINoMp2yxFqT
95w7nSjPL3rimg6KU6FPAs5Pras9PHJt+XAPOQKB8tVUAx3GP7su2LxZlM0wvPH7
/AEEnoRi51PAMVkhIt6+Zi6cIxAIkQHrPdEp++0w6iA5npE8i7kfFuzZXegAA+Ty
BG1+Ep0rPmfVPFI4dY6w25pjm7B/tid8Mg7nHskHQaGWEBQqlHAHd9XBJcNDMF0n
qFMLx9n4zKf9NnHhKVqehCn0YhQ/96wEg9pyKR+rpODcVMmFPa5kyQsVlqiCI7VN
V1jykhQO8auSPyLCHSRzMQ2FbzmCd8IoGp7tlNswxFFmMKihSVMJlyOVRUKnpBrH
Izj9fsovA7jaPLRdDjwyesRQo7v4vqkKyqheNNNYfJ0=
`protect END_PROTECTED
