`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ATEpmO8ETwEiTzm5b2k2p4sU30LGTty3TsOLoPYYXvxFYvnLrq1W7dth7RZIrmq9
QROZh7O/tTXm/F57IGZu2KWwm+gAIDyh9VltzBwl1q3OLha5ABO6qq08rHb670LG
eccLZ/GOa1dhxZksEE3kASA54O9fjWW1hLDNUVDOLLlM6w92M3Jq2d/rsuZBpyj9
soofE4MtV7fB+ch4qdgp/wTSK3ALMLVI4G+R2Oa07ploJcqAu694MoHQ9DcBNTl4
8mLeomj1T0CET8umXVugjylsIEvQD8KvuohH1IAIeerWAirVeVbBcwfsDu5TIt8/
ZWeUo7S4iFPNj/TsZT8utr5IzdMcoeryVLxGl3iKyRYSB7nFJKqx4xG48KBed2oH
8uBuhJMj5yI2Te+G27MG6lohRqo1unnaKuGkyUXYucQBI6E8GNyi/YW9P6QT22E7
0I8F/UconEN+tgYDXxmmgiaeYRNgnBozyvAJjwP6xdtDh5JgbfOsvGwxNHadIaO4
EQur7l9jEInIZYpWQBQWQOxbT0zMChBwvVio465zh+9AtfNIgfzffzRfOPN/phom
HQWfF5EBc6klgMEbj3BhOxRvpEqWFw+QKrkW5voKOMaqa+4mdLxF6ptORfO3sE2x
zPYkNoYDhCRTb0+8pjinNJlDSa9umUjHLew0Z7Z7rrHv8xJ0uNzZQmnn4QZE2Mf2
uCA1kqUP9IB8LCykm4o9D4jsnxELoiV1lszXoeb+1JJncVvTCqlzXZnTTvDP+Kix
MI026fKPPr826578M4DMNxFYN/vkIg/tplMitT5fjDW8N9g9wWONJPlbmvCXTuSy
iWPHgHKBqMIRnswk+Qk68v7XQtu0PwtAiZA6/sjBQZRAkSFxWyRymy5mTJeh5Gvb
3CuWDv3up0DIKqO6QR4FAXmm7/ZrnKhJ5Z4nh7OphlA=
`protect END_PROTECTED
