`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I8j3Q0FEjp0IKIBk0tnf9bRhZj2b6CMaH3naA8nYYBowC/vfGmKK0jyQWVjAqUox
Kdoqpazr6KcZ0EufB/D4FF8zvgdRn4DG+reNXjf9JE+jMcRhNhyXoldyB89GQf6C
yqkGGEHZ1faV+wdduz6oAdpfxdzBbjgfCTkqAW3F3gbW/INPmLOrBwW0KDFDFpoc
qfE58kaj0B86sFsJyHPvI3uxSZw18RyvCJKwTre/05ao6++OPXZtDnKqizbDwRAq
m7cICdU/iLMJptAYg+h1RTjrkm24aTkPzJzyNCY58wNNOp6nBmqlYvJXt13+X4Fc
WbB+IhonfEedFvQtHwBkf+Lx/9o/mmhDztHObFzk2xOxW5llgUtPYn2s8SU1+4nE
5HEdHalMM7jjUVHp8z8wuW8v1z3OOZjgNmDfehmtYZQxs4lZhBKS8Wju01Wzr01X
wtdsrIX2SDyEbfUhPpuHYw+8fLKyc6kjEkwI7NP8YQe2k+Pn860ctAyM8d0AReKR
nEmjR+fdniASNtLek7cdxCBnQdWpuZ3rSNDdB8biK4YL7sEMst9YBjyjWWRgHa75
EEAr9qio/W2FaBkjFE1i6bEJgDxjWjHIAZmfRzp1iJwBadz96NWmdRFXGsxtzcmQ
WaTJ5WyxnlXFGMkGabF3dLAdt8sfINAvsmwhowhPh1gtIeCWNf3/1a/6CL2Ovzm0
T/B6b2nw3650EVFTi+Yh+lV1ncPFZqZMrhP2N38Dd1z+HyhMgrHTCem7ILBmdrwu
O62R2lOfmKg5EJ+8SNSv0zJvXRzbHz/7K653xUiMsSwYq6QLqHDd7oYbeMQ7PgMX
S+lt1qKdMMllfsI0V5qXJ9eGOHx7os+MBInZw78B3y8EVP/MS1g6rLDZ9m+L6q7Z
snVqXP5MAu1eQOQ6l41T74sDxkAOx/ZM7wkqqsY8ewY0+sy8JJbbnKCQ3Uhz89Ho
IZeXACcA1PYX8qHYWOtX4KebwRZhS5ZycpW0nb/wIVfYuabaCK/bMFaRH/cvAZv+
VQJ9ujVk82V2DL48A7dJGtfL6Gk4qfkZy+Cf8A0LmH1ZT+KrC5iDNwAcBgCXjT/Q
fD69+MC32DRUds3eayyA5QGQs+6LDJRc17BjrjI+KUlwGUmugFbblAk15iNN4i3R
HzR3ItvT6pAAi13jtAWJQYtkyCu0mFyUfRZ0jhqggWYoz0igz2xnwmywsvJoWl+V
2SwHoFsa12AUWGvvrwVJZv7NmpUYyKLlqFDBIhtL1rZ9LSKAHXt40dHCbxVXKF7q
sIGXIpdW1tzJDmJPfx/GR/fioaFr/C2YEHt3zI6Zyb0=
`protect END_PROTECTED
