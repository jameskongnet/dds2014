`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vu2QxRx0IFt7mNbhMZMRRY4LR91yHl0exZ9yRNzZPPzUGbizgEW6n4xzz/Nj+KLA
09PK8dHO/Tm2egzOA9QC/RnCFG6xr20v3hfJzfrTPKZkupSMUKlo8QJsaIi4AuFY
/mjzosQ6TbZlfhTcOsp34ImZc4mOr5LyVma7VuQ1mgnQttVhAxzJ3B86vKVpPlXF
0kO7Dq6oHrfnfuFJiD5mjxPX7Hp/samVExS3KNMDfDsUzce5TS6MaTWfCh47Qplh
BmeszABNRVVzhhPpV2SMBG8YvZOAdO2tV1LEDiOz4vzzqBQm0zTrXFrSZTEREAIC
Rrq3zffAMwTTMcATCdzGfxdSRIbjTq8MW7B8uXYcbSTbMc+SAUtXfCPbdaIgi6ag
t++f+proMJg/8PhRuIeADJTHg+Ks3cCfqf43tKR3y8ZeZwv6q16wr0iuk0IDTxFc
cf2SZQ0QDAMa+UHgMAJM84NrGxo/KCM0121icowaCiHbyYcdlgFAeJv84NzxCL2o
xfSIR9uBhti32+a5BjLmnVU56vOkWer3sq7EWTzK7hJ98UvVyA8h8JyoVF36gbVL
Iu5LpWPZEepweoEIhJmruvtCbpzpqQLJFBtrNKFDrYyVnr/oKcBDx40IlO1c3b4q
3UAPwP2D8dNTh7rT0p2Mt/Q2TW9kPhD60JjjSHSBFHEzthfB+KD6leNMv1jj4eyy
94eEiZtxUCbDIpZKIVzcwMnOuyBi8cCiwhc+xBpMBOyn1u8d4nT83hxNesDU3HeE
1GevuxMYqDkOQcAegIRzoza426fDSxiTVHpdtS6Mg5MzoO/VAD7aRrf6tgq4MVPM
NCg2T4ro93xHdZvV3gCD4FqC9Nm76MOaFHRIPESV6NOU4heHWTPhIs5R3LNO8yJ2
e0aHs7jJ5a5y6OsuVcs4lBIgBYZiiqvY/6OKPNsOg/Dq/V2mvRmnkl6ov1nKx6fJ
4L/5TT4cnlITf2DaqEG2CDaZskv5hRMjKsSIXBaeVd3hdxC96HAPOzuvzimIjXeT
lZmRGaVAvza28giyMmKaxtMVYeS6zPQysY6igYt0VwXLF06nc4eTPOD/UFLOMq1m
cHtln/2bf1UkBwDOorQxMiPQXA+cFDFXJZjQ8k8hBbk=
`protect END_PROTECTED
