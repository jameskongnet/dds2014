`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oKQMgwPpyd0ye473BK7z8lFr8gsEtKQJcd5tzFkjhV4pD2V96Pedye+hzWxjp2gL
rpdAKBcvBuh9uZpliDZvCbcz+rad4bW891stDBaYYyDGBQSfpoLkdMPhjoJetfye
VhzfkkzkusY2PmkdI30lp7DiXDA3dAuvR1qMQ3i0uaJi6iP7Jzpb59eh72VCnqpK
TkXL/ldTjpWvzdch4fLdhE8rTF9vHL73JB+LmZipkpshfn8hCbmqF7O0R/yPGJjS
e220P9LQbKf7TIpjgwowqJsmvAvDz6X3+5ZgoWhS7Ev3izlDa8us8nQhCJpTqgs3
lKhcPUod0SjxxMdaEyr2cxXMq0jhNRQ9bl8bWjK7AV0UiOaYHLth1FfmE/6TDP+j
4L6XowNHs7tHFUMOgZqDe95u8+y/sbjf4psnCaLNX5XxFL3bTVfSzThZFSwjqYSr
j4aZ/7jU4FxmXHPui4rKrd5RhZpWjivHPj3tLAfWfEjdMFary5u/VaVw+CM1+Ai7
Ek+g73A1O6H77D9VJRhzwU/x6lgIJLNmZcpNVyThgiCEzUTHLwNV6BlMLnx+3v2y
g8Jk368aJhMwvEXsJ6rSeIXVKZjU2uynLfqTTFwGMV1mDyOKv11/JWAYjZ4Z/s7y
xePt2cimcV2OQZTbHLqCDVJVK/c9gGwuFd0tyXV6mLq+yaDiG4S8WhSy1XWnzgqM
6wb/1Y/z2BqcrcLLq05QpHUhMyECoqZuHzguxoImXXd5SUkpXm6iexoQY+M5lc7X
MwLcHIfbcOPjXM2kBLQsoNfbClAoqzUnus/JYFnMwX4z2oxH28qc5zjjT2dUCN2l
qQBqyU8hAzOZ6JHYxG/80K4YDwX7b7wmM/mjTFX8TLQppTE7719CagDmkZhzrLdd
Q6RvnIw4JwEBL+ADOA7cgPdU02n220TBdpwZHe5fhtCkg30cuV0SuRIUSU1NGYGr
8dQaFU5albkibdXr/TVKC+gHO3b4XWCF8xq7oq/nJoBD3sB0P3FhXYf7YlcMwssC
DEs34XOPeGFgYt+d5Pa64Tu26r6DbZHvfqeyytZX7MHVcpug4xPjsMVOz8XteNQN
Cn+jN2+11yeJiGdYT/UmMRSZVJOpXjjarHO/Wnf9gkcrk7XyUxCY+83IJyE3LG1F
f1nqQ+T0hOf4J+ZhRHHCzhmqav6f3AkpHcnjYqGa7dJsbHY82VKbel7bVxQHw7dG
c+QIr937UWtP5Y1WLV9jywwWgLy43zetu26OC4wkHX1P82ieUDAtm+8dbpf2fTly
qdNeXUZ8zfvceGJxwFxpTKg+7YEf9aomN9Y53j8i6ee9Suysw7RnR+9JE3NB+KSF
7buzaji/yJQBe1kGFDITCe6GyU1B5y80EAxfn3nkssV2YlBDCR6/G/JcjsHeJBek
JyxkCeeP8EXmxW7tmIer9DxBUdKSb51H/a/nmAq+3uui1ERcSPo+lWzRapvxToZh
9ndLEflQ33w38kaSOdxPPhw5DgTqCFEpZYUgpUsDrxXCtCEzAzMncYAnasYZdkxu
pzbSMt7GyT4Ee/26yvu7IKJ7YC9Fx22b2RZ3Q4sx5KIaI0tPaodMohZ+tmVfwG5j
AXaOq3+/wAhNqjAw320vIAQz20sRwNrdVRB/mYMaXsoXTI0GY92ilA0YBz0fS5zz
AI9u97Z8evbOOEEh57WelcxbwdJnEDU4RBjZZGDIl9jQQQKlh8izjpgk/Gp3Gflr
wqxt2JG+dB1AugI9z9qLN2319Oshgd5uXGOcK4vgyWUBF69DtvJxhPwtnaH9UALw
wa/vfnkJU41uCyYGs+1n+9C9Kkh8DDiG1glgcyeYPvBw+DRU83QJLTrhlDcEFM8x
jWVRkyUrjbDfjtXuj8+B3DIIaEJI+oI8InmFvKBePsYbINCcuavbyvBkEG3T60R+
KHWa44Nlq1xCepV/gHMgnvI42/mCnkLN9vhr6pn1EIhrjbxqDX8AdgDIuyXvNRjE
R1+41EJLL2x4g/70fvBUTBMn6RLJ6x7oXzMqN+w35AshloJMT/oKJQGUjqZDTLDh
R9ioc9ABGTZhYGajtuCQ39O9qdUT/2R1XmEBnY1A+4OTnDic/JRi7a/PADp2im6D
ZylgAcy1Xjb+jqyP0YOROnipjtkKWOiOuB9hPxeCT/bhi8Rv69qxB7IGAWkIR1Fx
gdeC50HWtqG7AwoiCOeAvHSGzLv8WGdCl6OdDQQuUaSgzYeQJZ++uCGzCaPvjbf9
PvciyZxkfrW8h9eLZB+q8EITBKfjLQHFBtTFci4cx0GVnLw531dnQXDpQL7hvhKY
WhR+RH1iiWCDVDAfUNELEe4QiOqEGVmho9kINzX2w9/OYsIEZCUZTbFVHOsT3zXC
oxJgxz6uj5ssWV/M4vPbnVnZz9N6UBOZPTZ0sHknceB/AN9xUEJbx6mCa8uNMOiA
fVa9PdDXeqXfYFAhuhMoD53oXIscIUMMlrD16MWvJMPBwWiX/LslnNKyXL5nWX5L
TWHa3OhNtLUmfikwg5A4lJiAqtTb5WjNbQUN9VoWrrln7zh1I0om0DpF602ChsAr
fRKYpopDZ/yJ6Ux9/Zu4eOHnk9CSJ77K5A3nlNZw60kCwXliBpzRxODZJzRAxCOc
vFtFmChVq2I24686w6rA4sTEzdyj5W9SgiUUMlVu99CHsVMuoB5wiDmH292FLg0P
wlkxSqsuJU1PU25gsj4wGZ7M+2dnmwznx4a9zpe6zLDQBDnrMz9YXQiftlfNf2KC
WIJXOEsqhBj4niGUdVyNU2Oq3YNeqT+PRLm+Lx66nRy+WcBimjzM08E35518JrUJ
2erT2hsceePqGfXKHGA/5RvWrlS456SAsTuLD6KLnugxGiVjADvfy+p0wWSZPrmo
AcSl0pDy1CCoPA7QdSt+3qF0RO6zFi+4aRVVZNvK7aws7/A2g8q4L9vDPqlq8M0E
iYyOgIpCVliXNCOhi5j+W8L0Zupqk2OjmCN84UtjP/4P91J/2V97MfGXt5pW9/dn
/Q/piXuq/vIJ9lH7EE381Nh/yx1tJmnNqKJG/wH/vcO8MiPJv7wxOyF8+s8SuBRJ
3iPw68TpqKDIYeVpOwyPy/xene4xUOy/Y87sLJGmzby6WKcmvSpqI4eUzDtz8p3W
9Y6+/gP1zUvnTBg6Jm2M/pr5gF6uBBTcGYoekx1Ah18Nivw0FTKWFUcoOaNK7b8v
/DnW/mWlEbdHJVEn8OVFzGkTY112OLURGxljplcAdaN7xyGLKiJ2jZUf7qc7ztqQ
1ob96lmlmGp9/XFe/lRHnJPkGcOijNe/9NBrhqipvlwIGV6fEhxDDR8IqqsWvy/A
+eI8xfGpa+iH5YJoeM5oaABlsIjIeTe045JrwCS3LxMKxiEdtYzhG5Az+u8vpysj
VvxMrYKmeQqxB0WWFlzArRjbGR5z0oRWZsPm3ZomgqNQ4nprI07PkjC56nPLX5C+
nLj75wWY9wmDRu2gKTAcAOkfw/D9OlDCMDJAOwtzBhNMrONgHxscBQjmrIpW9vxw
+ud7YxRvzviXBiQpRD60H+dzUnZUJ/1zNzka44SU2g2fAtVsPqLjSyiqcXr+olpM
2ICghVtSqWZRGTNHiO61jGVvMCSp6pXl82xe/cB3h9/q54MOnIAHEkVR3c8yVEEk
qG5ScOg+LYkEqjXdbxLRRDhR39xLWhw2NElu3uZKmP12rdPNE1bLy5+9SjNzPKIt
JqP0wq4QmGyK0Xbe3lxVrBRhWIWsxqFKRXyxQNPcs9Fnii3sFypC6UXjyM5rkSKq
YCQ8ImqsbRYsCGr6ll3pwk07i1R9C239ZYm6l+NFUdKpkcC9rJeFPpzYqNnYBkW1
KCuZFKNFTTAXb1S/UwZY+9XGsm7dtaonFAVh/zh7bkQQso5x85gryU2E9CbdZA/I
rA6ayFhaGLOZrr5PBhSOFkv4sc5ezrIDSYVa6re7TkejaoCW3oxnOEXiGPhFJZAd
eAUWnElHjX76sQjvC0vVqoRl+6aMrWYm9PLmWx4LSwjJZ1C0gFZZ3k1/V/2/tCrp
fjFxxQFkBcx9UI783pW5QuFAPPPbsZFY8uFKPy9oQNhw9IRmQFKl5l6et7W8/Cxw
CrPzvZPg9tQe1hi7/aAGXO32VDExn49PUAk9VgGhU7P2EPBSRJzsfG6A2xtot/cy
AcoGrKZeUTbTtTN+JLOQF4RTS0NV06bHePS7q43AiiQSVRScXh281KoRyjwEyZAn
f3H3T1X1Ef02ZT/0iPMMpVkDvFGs9O18OHNVFhwsmW7nuekzlKwhI/PWohJMjqqc
HbTHOVW+O/NShX7YyNYAHdZ0uDkRFcmUfTP/4dz4spjIN5ovdDqOXE1FsUyqLS8W
cbQHm4OsTUrXlelD44SC0yctpZu9iBPJ6eevPEKkevJFp6nG1oLEg/lC8Cw5nG+m
eYzUFdUlQE3ry0syAWgUJh/RNJfJ05DkRP4cSUhRaQYY0MobME9Znf4vKXzUg1+3
zPFeQP+x7t+Y+2o14HKfxn68jtpVqmPvj2Ta0zFaN5ef8py8enyzNRmo9tkvnNwy
HTua9z+PXp0vdkJdZSWAzPWJqBUlxtweoIgBOOq64zS0UU/hfyAUzIoJSezp8ZN1
X6gSqxkkyfJJ0/RR/8h1tPAwpTJPFGzPCZUa6ywVOU76sr9cRNSPYRs51Qq+BAST
b+W2jbKZwi/6meUsin1ovPDU6lMOGsU/b88y2BYe7omwG6qDPLgM9zhppXUISMLW
ez1pWFnn6YFH5PIsEzQ2IEd0UobzBkffha+QTUdvRJhaOCHZGAjZM9QyeeX2gM6j
414s+EB7pATo0k2ncZIdQtIdyw/LpGhTLHI3zH9L6aRU6bd6Pxtd0TrNL+DqnlM3
iSwJh3kubaMX0Om7Q1zSME5hga8/K8m+QdnvnXLRcL4S412tlh0Sv5W0sECtdqWn
nG4GxMH9011d3xR7d/D/hHtJ5VjYqiutkulV0NFYnYxCqGRYiYxBEflX3ytohGj0
RkBeZVBHYh2zc0ekolEtE0BbUA/hQkBw+ZOYmYIyZCRitNFxhAPnqHh79mq8BLQQ
OxuPW+iRMkCAGVu7tWe2manbQVQ3gd6ZAphFBprYjJ41TkErEQyXl3F/jLcbAb39
Pp/qmHKctevz28HrIjr3ebZr23RiOVmomEpOA3pYDmoabTFD0OCzKR40yYPMogT9
WGdt1R3mdp2DGGlcfoTxahlGZfrGuaN+uqudQ4qt8FEBazJB0WKyuStqEa1JQx76
1pPxapLS5MoWPaOMLN+aybfyTLytWqgtPQ9Cful14KFfKVSeMALPJSoOty1zARdw
+EpF8QLcUJiHE4HGMMKh2AmdzsF14boUHAxjVILvkWjbY6tpt85F7ElllfiEsUlZ
K4OJwFulxLocGlmqz5K0KDv1FxcA/7HGrWPCjGk7GkVc5u1V1s+V3UmqT6qt0gZ6
IToIXyk6fNz1Qjlswsoj377ZjxYOC9rwoc+a9SgI68UNAmmqyGJbt5+sEE0s2c2w
yeaxTLOVnFGB1QWpQbUiHEUMbKUoetELcGV152ieNNR+7F3iwSE+vm9U6Tm8yaUh
XZ+/8dknrVTrznAjUuWr78D9ZzeFI1hvDOdhteA0QllIF3q1F2IbxLnZXBKTdEUB
MfKRrhxugRu/E0g+yiBasGEKZXfcRFj1K50PkdCAgVcP7J+Rbh7ZWLIAhRa5qBgb
WefB4yQnFhTByL5R2FAmgPuRD1BsUkiDD5Od4CoVrIm0faUXbDj4QtX9BIHl+IhY
l2ZL7VDcU9YcsEvCIh3jmDp+McqaodIwYIZXyZhlYR9m/H22O/8SZ2Z+Yk0hzvvf
xYA/khPwGXh6OXJhSVZ0+adI9noMcWi7U2teufedSljx0bEo6hCK1lqE/jJdCKxJ
jvMAqkhfp1/CbzJaYCditt5w4JmAB8I0QVBGF5YMfzQTe2l5yHAZmEmnevG+skQU
h+ot91xGi7b1wa3SFoKZejgp6ICzvKBoCtR55RZ/LRqk9n5S1QMrMtSO6O4FTJ0Z
7853+sSPvrCNGSW5gyRe6O0aCFvOYiYFUtjAH7NJdByKNbjchF6EBZeiOBlDEa4w
/Tnlalt8NzJzJbh7SPhOBDQzM4qHRvtmjkSQskOk8e1gIqMn4Xogl+q29//neFYY
zULtoAq4FPNxMVupPuj4gvqYlYJQkPMRGoGovplKWj4kMPBYRUDU9lNmW+ta45QC
q7tGmsYBJH0/c7y2pwYsPLxPwQoW4TcLbjQM1QJTdX9pOnPanKg51pDEQ3FZsKtM
k76NrJZ/QmVHlKUgNpVyuONLyp9BYs3KSeo7onmh7aGyt3O+XoiVc658gmzLyw61
0ugwZMO6gMHQiEqlUmfz6IEkrVVQCVBlB5e3QFlWHNAxbTiD2oY6mLq6vL4n19Ck
MT8Upch5EPtHb5yXku/07ciP6gQ6XPblAZ815FE2bZ/GhKAG7QJzI88L8gZQk2Io
xWiII7mue4tvTLGgy9ZQgvyXkmYisTCBIeH6WHCG8ewPeN2PaYwYaicYT4gFS/rB
JMdW7s8gZ1mBGb4p3dL5OZKX8vQfTDudFCiSxIXH7t5VPWIlUnpjMgAU7Y8m7+Qh
OMjkTO602dvbWV6HZQ6HzmRKU3nNTIEHAZwpMcnBQwSUdOh9DGzbFKsfrf1jp8BH
NOENS+yLp9uctsjnweG2jLrvr9EQFUOq6hUe2hiUoiE6mWRT00cMP6VCLVsIpSsn
ctNNTHC9+pbYOSeroueDHLqpQlKbl61j/OMtcmhQTlw2j5tdnB07QsiCEgqDHoBs
6R0Mnz2Bvkg+Vnl/qkmznCRp1rDbtaXiLzKWCssQiCk0pQTFpRAOJ3Pn3msGlb2B
GsH+Fx5ead5rZgJwIHqyWRwIoXbt7D+Zfyz1cfl7JL8dX3a9+RXanwoPbrAscnYE
epNgno9y28j19ZO/Egpr0Orh1LguycNjfy5HRhgctxVuQcIHgSmiSdT0xhnyvdDH
vfD6mTKpGJtbr27SRgoxqXd57yIR2xdqdqeeMHmK9p0wzRdXhShiVUwexUFeLk2v
FdOzEzLiYP/HeGV9N366MTTBJdxCbnQouDYkwjM6BbHJYrEqpqnRFUWdoPMfnpM+
igyTsxGhHsjV92DTOsUNLSVH6QUbZHeJkphfsTMqKKpRM3roZGAyU88CfGQ4yd3R
MjRPO2kSABX73B3tN3vJld08LtHUwY/7GVmt3mks2GMoRBfEYdt6B8Abknx2YawY
nQ1UoV6lK/1r8LOFC5Yq+T16LLJLRI77RdRBQsr2XCRNYFJeZey05kZF3eDK2uK5
GSGSOwJeJkmtT75HClPAYRy13BauSBiR1ts7s/Ys78vwrrVZGZiOIayVPcuGLuVq
HtCGtCZKBa0gxbXIxlBiL9M4sVgjo1htIHM6v2S358BHKXmVT2hejXkjseaElzP1
Zd2StMJ+sIPQWeBkYla4CAQ6myRST/IrNw234lo6mgpqAm5pF24/O7865xHBMOdU
1OiKqCaPBA6Svc/HB01nv5lyCqjc2k1UE4nKbFWPBeJelqAi6JGdzzlGKHGqeg84
T6XUozdqacgMnnI0DvJM4Rc1k6X3gz8Y3oVbVzhWn6GnetdGGtWy0Ld+29v9X/IQ
BhkBiml3dPH2BXGzIvcrIT0goQSoeb9IrgZHGUYsQIPiEsbx4A2RJs5A+HWmgbCT
MK7ABqiU87JsKTj31e2M7hMbGEKi8k/mQbLt74jEdYSb3sQ0x6Joa3K8sPP/3ugA
MlWzPjbYbZ00UVNR/6bqFKwuc4qcaCNFbaF0TPIVc40C2CBFvdqL8fJNA1RbNwEU
wzxSJpn0tKEdZNg572JYUmbZeTpLfGLIY9Ru6zBQM6n7fapDnY2IudZrylN/srg0
7A0yTpA5QWm0z2BNkBuwJOFRYT0JBH8X+VglVcXRVNFHsoUKfFLDk1sHsXpbUq+b
Uw5gdFvgkF8KqScXWZRiWD8+vdIRI1PTgLj6NShlESnvHcJuJpUl0VKze1G310dp
XSRLbY10dhCajEAgGIV2VL8KLwle6WRCIdYrzSNcVdrAi02JHpCEER+AMVQ/hmfJ
Jkjk34v0NtW8Z3/qyIeBvNU6XfewyHH4PSeaAo3JwRcXOHUGzGnxswF5Fi7reXvL
SIsGI8W3whiew14n8jpC7H8QP5JuusqKz80iA2t9R2m7BlbeS674zSwbn3kbt0az
i5p0+kw6hI/th/y2M2CKO72pbRfFXm3M89cBtd9rMfq/MkBpRdVRaD+t3AdogO1V
uxPUWL8lbzeHIfEJPBhim0bGv9L/d7p4W7+SMmzQTBMD2NxdXn3SMGDxffbKIvC4
4T/Y4ejavtLI+9zvfaiD42RNwjDyM8cZsxeeXT3dwRJR1SCpo5FFA53AZ1nOa3/B
hT/DI4WfzmMpftEkS5TE5N4I+9s5gyvzIOuGLgpttkz7UAMy3Fu8Z1AUVKp3fgrb
+jCILexN8/zJ5u1P+MA+Nz30043lkHU6cf6r7m8zZbRzVKxNldcJHAIO71cpBrYQ
ARDW4vjP9fAKudGIzGAK+UxG1WtdAyrBKi+NIh05ldIKesWgOHP+lGc0aY0hC5gE
7BGucOtGJMudgY0EE9npzz6fjHTZzPn8Kc2fovObpIM5y0JGISmpL99p0nUXA7/j
pkvUjneKlNswGBdCYuAKqdUcrbbzaQjUfoYnvcrZCqgZgz3zrnhgl71Ft2b53IMn
7lHVM9hca1HqpiNFYGjFE7ga9WB3lJ9b+r3jTmMiipx2Imao8TSfbbYc+yfquEUf
oJROzRK8sBLGNW31X7LBqxAV375VhpymyQlsuDpaalnUT4kTVEWXZZruODc+LME7
emVxn1YIJYM3LuoMvUNwMhiNX16EH9M80DDNrq4PIm6eQkkSwaB4k1j84LbYBj8X
U56Ow1d2a6Qdeh853C8ifZvSRR+zqoXl5UfkeZE4DOO1db7bp7TAGnGV+GYic4he
r/EaocQk0AX+kvf3T/uSJcqyF4xfmzL4vThXnZ5Quy2p0k5Gr/gdGUlReMvHh7nO
fVtVkHauu0IqH7H6droaH5fYwaPobTr0blE/V/7ZjXU9Ciq0MjC8V2UL2PQ0d30o
BIy0tG58ZXtgVXCO0GJplOu+qbsibKtHbxiFSioFDZHVSxMB1A7hEPQSbdDbpR61
dJ+F7Uc8LtmF8XIxSwRZtjK3tMORtaqW0XA3oMWFaPxf+Y4KqV2Qd29C6nxOKi73
KoDT2f4rerV41DlXl1uIpLnVWcx0NhXEvfTexB9li/KJezXRbBO/JWBf0IBMHvqm
/+Tqjn9l5pB4FO8sHWdEuqTU++Jlc1mmENB40hqC3Ys=
`protect END_PROTECTED
