`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ffznbvZiCeSq8Wc2tZJgEt64a/lU+fm4tCHe31AYWK0JJiYtppbBwkMbOAFfDpNj
7RqGK6TVpe44cRGnHrNdvRuFfGhUfSCCzJqQSEh/7MGYOOK7cOrmePzhDBPRVJJC
vAE6Sx3KzDwwA5aKmQbd5SZFhUZ0cx5vaNKKSLIgPGmtLhJUIuse5RDrM0RNInhx
/DRDMwR+Cx6+leZynPP1sjolWihzeLuk2/NjWQ1Dc5HSpHgLKhmQrq+AXZr85ivR
Tisohw8pEKoAt7++tFzf34hFOrZMGlWwLz5LFdvN5wRIEEOObqVgWqAJeM2Vow7/
aFgtKJM/nDHGOJUCk1Aa/415gV+QXMX6wBQpd5GXJfccoFoJw4BnZKOJdcHy/fR6
gCrTXrsy8NOswz5GRNmxeUtGz/HkPheOhQEIgzlE6SHd3dxSvEvFlfsA9tUtbvpy
vL9xJXWmfLNbovqoZQpNzCLBJRUTEI53724C0QBQxBsR03EM9Zk+/ZtFntFgoYYo
8THwJdaDmZDjD09lRxP9y6VW/A6DO6CQI4fLGgupndH58HiOCswmSD4WvKEzYG14
IH/YP6VLBr3/LzxuR6DhJ5uCa0+qJ2BmAlfVhBF7HLjx55i2Gw5TyBjIXplTGrcQ
OU7dznUoiZ+1nTZre2GZDsTj4fcku3/xPWojIRHqxyqpOrqb9GLjgzo1Zycs70OL
3JxnJE/oMfnfb+cwdtK/3C2Zphi09B3enneAVvi3OCp/5oooEuAXzT8pcUbS5fiG
xXlut9mMMN5jtXqDuHEbMLfgeMr8AcMdqF1LzskrNgWPcv4jgwCaeat6UywfHHda
HO6ov4RYrFRrW7HNwcgbI0H+3rzKOGl+42uMGujC/YA97Xj8q2mMayjgXzq9o4Ut
IfI+CYYBBh6vZQQUd3PoydSChzfRvc93hWVqr9o7au4PwCz2Q27Vb5xYL98R7WwJ
PkxLhSfcVA4+3wj2lP0yiMG5U1kzkxMxZcpEXDvJAKvA1qcdfT1Up82gs4Dk8XL5
JM6Q8yTREMzJeu4FI6x4f/TbgcBdI4k8xpPu+b60F39GglCGHYAsG0C7lLiMDTdf
jwCcKKHW47Nr16yE3A0mBUiG/Bl3AsxdEIPLv0ixioDgFpUBcQbRTkWX7/qNhkc4
NpSP+gp01qtyMwZPAz5ybRJ8dE0Mv0DRw5Ml5O08euN5hvXEGnvwOE8lNumZFrGa
JLWp64yzzZcbAcxhdzYDOemETkJEzS/PKQzx+AdI7Zld8hC4B0YBtwM6WF6XsfoY
marwaOVWB1mCO11Qr9TyZz03udYTKqOjHEFstjNpDAxLa/FRsG76iVLNm2zdk3vg
xSgg7FsNyzqSuajOEHc+tdoCBG1sG8uT1GG5nYN0umlAMvymV7KRiILQwtDahilB
M+PqwA154EpIxwzwT6gB1yrpUakkpxfal0f4cjSQXCvRC06LFGaK8UYD+oB7Rqpt
Lo44Xuf1gcfenrPp89fb0Q==
`protect END_PROTECTED
