`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dr0Gnb71mMWKGY5T8T6ayjh/+vPnNMI8vB+o1MxmuiYXQze2/56XW99om4DP7NoT
g8TeuglT41YHAE5CLL2XnnLnKzwoRsSXrsgNbHWmwCER6zePJmp4A6UehqqCMEuM
bwuFBJRgBPzfsnT0d9fIHHhMxn3lq/jhWEwcjknUZxZIgKHmyvnoEs/EWZHvzeus
fgNeFBwIa4TW7D7xABATXFeyHs9Hp0KU4M6O1GtlY6obw7pkEH+XvIRUdY9RHEMe
U9uJlkbDo87wMb6355g1DbuaekxYBAndcuccHR4zUDu2tpAmPgG1AvovWiu/GyaR
U1aRgYIYkHBaM3xhJGR+hoELOMPxAR7523yu3d7kht87TvWEOEMSfcZuvlcSZTHF
DAaSePpsSm0ZSF/jsiWNTm0d7U0utCUtlCOGMMosQiK5UT8misf/zvs5dHY2Ggjq
CF/e0mA0c/0ipKAM36koIQD9pd8tP1wHazL55IT/XB1QxP/g9XLcwUKYOVJBgY4y
LksGFILNrBme07jtJeahJhAGKG86JmwgJ+7Hm+K7lQqdwFqV9g89TVIQ+yJBwI7i
N9qgrMY7D4zTA69/f3kvEc7CZGU3XBsXTfjS8r6S5KpJOcFeJyzfposTtTl5UPK9
58kmMjIbjpsts5Ks6OanjqgXcf6KGk0ZTDEDNzNsvLXi5twLTHZpsH0lVNoYVGdC
5ix3qB9egUc+n4qvObrRA1S++kPLeL+nhmxC6Gi9fS0yjE7BDdrdq92Yzne26Vnb
Ag9QQqrnWqmB37EEKJYl1cuBpODOxx11s7MfrJmbWq1wLHI9jq/jJBDys5Fje0My
pAjjsFuDY79iSZQTGvPzfF0zAqvgYz1f4FPqPQDp5Nl1fENn0bKCoqT9EFRIMGg6
Jebw8b3OnRvTYKL6VDo3zFD2chmXKBj4wlt6WRcbT9NvTThL97n5CA2e5bs8DIcH
ivl2E7jbg7tQnLqt5xIwBDFgH3GFX440ZpIdjtFwfRNY63Smonb4JxS65H+rOJSP
1x7PUolz2oafeRFF7S5niiIkxS9FmlVt08HJWW03ShOeDEWowt6phSIyc+ogx/TZ
w67EL1HzozLXPD0grKt9qYozReMnVy0b2kFwqlrStgwCjYl8bcqJuWapOFoPuXcE
pcWl1jSLxkssSR2+i8sdDI77N31HjQEHO3MYIsqpJNK5VRbpkcunVhgRyRWq1kzR
KszL6KEq07mjyA/9M1pjMVjAjR9M/6QqGQDYkr3UnGGS8g06kJiPiHffQHTCEVEW
UJb4B6TklB6nFmCZxSGzBCwRAPos1461/gruvp+TQHfWfQSaO45o7WUX/EMPDEkc
IXpxtqCymV5RfLnm0+O9X/Wom8bsscwKXDz22azho7K0qlYbjOYl7Zu42C0MEQbt
mzuPJdOyGtfUHElTgmvfFtQ+tcs3kJe7H0pZ1C20xyUzSc4tiej6Kr12whDxW29s
ecBFnRBi96L8v8+ALbv/2oP5POG/enIMGVlF9bWOIjlqZERezJ/sENMESfz0Lu4N
SjOF8+L1jmg0itzx/ixwU0OKFpYgNCGBhqudHlU2w5ZT7sYobPzz4YXfY28EIFXw
Dr8/AfAC7m1rnXXRQ96lGAaApmlesd9EkeIga2qIv5wT6zS47TsydW9QHF+a/WzT
Nk7HGPrJS6AagNlqkqH0kWjmBG7tqDJkMIqIVS0EhBQ1oD7YgJ1p+XK8waa/uESy
i2TYX+4HSgKF6QnK2wx+xmCDNTJbB35CNb0CreOT3E5iSDUugqobMPPbNKsuG1t8
D9Y+h81YyuEgyA1c+a470Km3cOjfHvRFUk9keVzTbi4yYDbIKGCYIXPZACQqHKBp
pXm4XZSxqmlavWAv9MgB39eOkaB/SFAnZ7dLpP7pCbIqJO4+euOJsNFNWGPsjUeo
ChNCfnvP6LxBKs+6iLVRRrhXgut++Jd8E2miu7vFnN2TNI7cE9Suaun7cmNc0tE3
LFi4TbZ8AWgi4ugkYgHzEtxunriEz/jk2HAbV7Elz1/zeUoqf/ZUt+wM/b8ozDL6
EHNVX5/J2OF22emkf9O7Rzz14DcmOkcYGaX93lphKnF8jtRLs93dHqUGcPFFXbtZ
ZkZpSqlTHJIsSU4IqL5rFo+vOM0wiY65T6ATl0YSK4wtXnpbGCxxD0v455D12MsO
kxZZDu9lH7oEiD4YmAhJ5Y9C3WK5YI8NR3Owx8i33ruo9lxJo9ppeOByezGjmnxp
pQ9qzQJ2JLar5rayIwNtbbaP8EU+865XX3LGcpM0uKwKH0jUArVhK5+ssFHb6P5e
6W9Juq3e+Xhz2Cc1IggTayRJlXiPkenqmunQuK5F4sqcuIIsvrx7wJe1xHH2W9G3
9Ar7KjVWGfzxTlM/a4aDbFgp45libjQDZM5JhPvSw+b1llp3fyB6fk2Wv5rj00wU
hlg65ARKTqJN5IM7ICq/nuwrBCJCAY1mYvFyx78nujL6DjEAtMmHJZAkYroeLW3C
dZQ0NZI4XWAmy/oPUeokXXEjmWTNxElAZ1puRcKvGrYu6Gb+FORxU5s5Bdh5L4Oy
rpZtl1Bv4R8eo+u/duusamv2YZWC2R5/742TQDAD2lrpVAIskYBYqMiDJ65azkdw
Jw2lPsdaLl4H/+/YDM5AEsl/aRy7C/mG7dNdL6HWsZx2hI0BY4dQxtsK/ixKImps
NF2emu3zOfpCUr6zgxxvFqjuZy5vmByiqrsGLDkm+QEJG9gGiZSMwDtNVA6g/Lxg
tjrRt8e4dAinEYBKuJy3+okoVlwrthyrFEcdoc2w4u6vUnUETJNHShuEf1EqkjSJ
KqRMljEOB5d61bgvPhpjnxtUz/F7NBwdlo0sfWajdi+DX9WclaYIv6+dmqFi5OKK
zimidrGyDFIid4rEw2bxuqv4DeMb26ba/CgCcr7koRdRMpf/Vc/rt+46IsTaDNyf
06zXOiaxP1tBhgjd122vOblOCDFD7IhxlRnoWyH8KBOcS6AIwqXP9l4iQRT0QFPM
qbuBP6M8G7hYwph5+5S1Xaufey1ACG+L7cVMNuttcFn2gRuVtqOvL9ASMGLU9MQ+
yXVayoCLrNw+ZTHvehqM6L/4xyyVAFNDBCM+iEfdpFgegETBP/3/M0DBeW/+hyq1
8VtQZROj1ZW1OOJoDvi4KhbF1DaVdCSuMsCsAoXQEPW0Y5sRTZUarZKyI+HzIoOb
795lAI7Wt3YTI0YtLoeSIQQR+o+n4tY+96dUzsah3A9utW441x7snXpBntCkSla2
rBKJVI6T9y+wjUoYQAgG9P/I9KSIuaYSVWKDakXqwXYbjBYV7inuW/Cj6mdmDbT2
YQ4ry7k3OMyQ8qDM7T2Endbjt0ljlrgkBCv6o4Xtnz4WZ8i24eb8O27QwolX0/jO
f4DL0Q71xChyJqDPE5n38lPTbXnCbgFPJdDxWB+dpBcFMpHy/LVVatDzN5Rer2V1
NXDzjR8pNAfWLV9bbsYOw8/AJpeQoz9wmsPEcKb/FlOBXRpA34LMtAaRHu1CM4Ev
V8PnTa/yRczH625MMR1yjDFphUYlGA/jcXMBwkF2iP/IjVfyFeX+zYor9iNWmeDd
eIBpmpP87WOOmLw4MUX/fEYKVD5s9bV6hh+kftrHU2KMmdQb2588Y3bbXQN6wkGn
uLaCOf6eVRJw6DmDWuWU3mlt7e37uyxyrNvcXUj8+LJpULCcu07clpN96z1HqT4Z
6qt1EwnDZNRGCj8rCBiFklJo8namgcqpfyrpAdax6f8NXRrR9v60boldhj41nW7m
JGo0tHQwyHzTaMh4eJcXaTV4COKO/Mfu6PFjeYomCcVpdzG46BIO6wREcjWO85ag
ae8ucVRFA8nMLcXJn0Vu+TSJ84mGkyEXEudZpegKuM2GEovO8s4c/+qdw3BiIBw3
gXXyo/ARStqci5/aq4l+icsebuzgeZx7CrM2nDLC2EtWvZ3EwB0MlsNDWrq/qjat
EsIZ/Ma1GjcDo9BEk0JlJF7tazHf3FqI7VMEIsvQTnsjLyHUpMPkre6pZ1vxMCe+
kqJAWKOiI3rreZwmDp9Bv6L7aIJB5stLaWQgUWe/Z3bVjjxKYyq+/mblbUDyGO50
cjGheYT4qMvvY/tJe2nceJaOBtKxjEq0jGQzyx+lDUCXR/uSShxqyJlC3So7e2HX
x5ImGf5a/20PMMv2BoCWizmnJbo8t/0GBeOFPAiIuz+oF5jBhc5P56Q+A+CdY+vy
owTyVOoZfI/2sM2yyfMlC10zD2GIiBBGqh3ZwbbBMtzz+oX+p22+FYHfi4tmexSk
T9p3xw6dub76a80yaLXzPTcbs93C+5dfU4hjpCT+OVdfpU9t3T2M1+ePr2e0YFxj
7VeFMYtO2i9H6qQ68UK4FC2wMMQ/ZevIJbcMobUH5d68nzv53dF1hWkuWpjpA+oS
zk5RdtnOnTNBXosp0itTca8TaICPCyg+2iFN9VIOs3X3PpNvEtAT0faAvQvfAvfO
EJGeYWMshwlG//7thcRoarHWEhfh+JRgEG4tFFmv8lg96fFTUgj8FfYRZjHI6sJu
QMfVB7C2ZwhoqjTPx1VzCbw18lVyvT5SeqCL+MzOoIR33RaOQy0cNB3bx8hlFEf2
8cgjJNaGTlFAQMnWhqKiLs2QVvpzxE4c85dEdeni3NrQtGeAVeViXnT8f6cnP6Nf
OvHimgcmNBQpux3qtWK4/BzPPv0hIJBft519ofxFTZyTdrW7iF91egErEIzgNn02
VbuBQe2DtL8xoJVM6zw96okkuCqhAW934QJvcFHmbKP+4c+b4DbXrKO08eKb5dto
I+EqZ7vd9w6BEfqfDAlJpmBrA0HEPX9FYd0GpNkXUwHY2+XDeCRMx9g0N6XDn3A7
zI1zz14RAh+U7ZehCYXYrRIIJvZRkT6r87NqC0DpQuaAsnr5bQ5NMPYUcPZH1U8j
+3rAp9czr2r6/EDp5fWQDiSy86AOqOT9NOnlHd5G0AgdGb//juwr1J9Jals9vB8P
brRZ+7QctGSuIe9TJl/4VZmstW3EaGlPY9SygXYJ947IgzUPnWyVuzEUfTMUN8E4
vI3o/9x/EhzU9RMGxpcW19Ac0+OztGVrZlVbQTATg40NFfcnk7zQiD6TUV17B3jf
CONP24bx1axGMwS3+pVjzmB9AVhlBn7BJWxCnUbuSySn9vKZyDo60VYnPugd4gqX
R5+pFXG0nkwmlDqvuQZ+ny/JRgN27IaYx9KVqa7qZ08V+5YO9Pf5WSd/Vz9/wJVF
VynMvybmnowHhAtGD5sjGkf5/9G23at9uUWQgFHa0sG7Yn3EAJPNjmHZ1umhL/1f
6VcoOfgzwXmu5YRPsW29EDj6cB/QVPwzh1bdiAZrVhljc/r71gcxlk0NUw+HXCjE
keKlVIKSXTbZwLXqhK0mMJFafeKz2h/BKoZS8uMDzPFO6L9oaeBKfjocUfdwP8I8
P6zHV8GQgPfuH1jv0HzvSJZEy43ERY1k0t9XxjknTSw8i0JvmXdxDuG5rf9v6nJN
ori8zqm4jdeQVBHh3qYsTJQjEz703/3o/ADWVwYbSwwndATnASnVSLAOOeIu6/lg
wxaN8dLKaooXnz6FHDb08XMd+Ykz3gt8Qg+Vp1TudBch3x8Wamh+kDVeMsNB1cVN
ng8z9YneaFks7vc7cw63ERQEocCcY5Rg8eQInAtnZ5JIzOA69bXe9Q1duz2Q1kr9
287QOFuE7vPuGrBNNX+9F6ksGIak47lUTLljv7zBTIUiiMuNeHYANHFMXeZDuzWz
VOHoRqLe1H0fBTokZVY+wk5nSHz4TM9XyrmimZKfPU7SAyjLQd03XhsWtjX+mRyk
Dc/zdHvvOQUExPj118yYPaXvVcaUU4AaAtpW72VAdCE6gHeXkMGW6139kS/OZIiM
K9vDdCyDvPP61oE1wYCS7hYDEU3NBykFdyv8HxjBEl/v7Qn/T6MdtyhXOzgrUBsZ
r9S6lxPcevagQ+cZnMNkJPe7PSL6Y6fnUfPwmJhtNdEo9Qr4oLCLqbRMDdKjeA6V
bdhUG0SPPbM9zVh593iyJKQxjMHzawmAXnYpMrFBFzQ6k/DPejJ1+n5Qa0osGi/3
9tWzGHq+lSvLB184KbVRZHr9BWI1K0xVImdxEFDWpe7k2oLgOO3cPW5J116yOuoJ
Q4XqGnyNEXsOcbAoOpSx4TbeBPqWj5kX/uCgZk67J42JkqmdplCGohMg/6+KCcj1
S8a4zguRNn6RpJu5Okx1Djp0z5nJhT1stvSkTTFd1a9ZN5nY/SFO0VLT7pPZcWep
TzRL33+6sLFmcrhxalXGpogUHnXgOJBe8kozsimgD+DWoFV+YwIGdHF8F+nRp7xO
2rzmlBf3Pv/nFcfzOm7iJxOXF8aQsZV4Svwou9pExpA8q8uxBxsXVpMpTSs6onbv
ZiQgwGP6uL8zBEZ9mY0rpnHKQdsXQnSn9xfot8zVQ5YjCvWaA15BAzx+M19tgm6Y
htbUAzZQhRERu71e+1iowWuUTrUyats0kWbbcPF9l33JOIxy8YapoBrK1aKzgV1K
+WxgtGS/4DJ/n/tj2MiYqebgV5YTVWlKMto2ylOBkwtJsBWO+i1Gw86PeONr5GSO
rC4aCuzBGpfLWefkdXFR0rq7tKKRyVKp+ld3U8dLh4ST3lZeFFobKybkGcJHwUXK
FEdFmxKrUSH7cJP9cUS9rjn5Hy2n48lo+Kb6K8BtrMdlGWgbjkydTuoZgL375Vk0
3R51erL1YSg5jjYG1noD1L3LuOExZUSlJyEUT4z1W9umA1c6hVG1AkXgaeK1gwEE
JmIV7io4IYT0ABIfctevUaPu3A3ef23yGR1dRoKAjYSAoUANhPGeDHK4mJjdcjCg
n6eoRrHg/LZquG28ETYAwTxGpj6Y3O4OkDGrseUgmWZKbrdmN+ltOLuneI6pl7Eo
PXeZaq9LMEyhrqgKqNoDBhU2w8SRbeBxw6gWtSQIueBFBHmL1ocHmRoMEVSNT03N
XA/Wt2cpgnrO0eNlpSUdCBTbkrpM2JAaFg5V1HnNmvqedjRLIBnLE24CPZ58WmOi
OasS45s+ZWN8ButbpgvtlhZTprxnIMHLvfLGP2OQPySC5I0wHQCsO/GNhqzW0xIm
TcxUEasYW39uqyHGbE8Ag8PfYYGPaug70DSwiDCt15n3rkRWTaMKNlr09utTfiGl
IhlEJaYd4zde8I2g8WWBcNgSGq67LnytPH0gDnxCA4UjVcDr5JOfq8SSQtQRLU8S
2EMTM1vJyzhtZm5DgiAxB98DqVhy8f2XouZKkuSwZE9S0E3TXaZMhQEZOZYGXcWS
pYD67B26/TGQvBMGi3zGDMkyDISj8N7Ff0MbwvLKc8ZkQIqj0WoGL6cGsK1AyXBL
TNLhlPT4YjEQL6iZkvxSNuALVGxdU8dLwNNzB7LFZId8BJXOMDJ8/HF8HNR6UxtR
Q+37HhmtuL5o9TnyygJqxexyAhajDBK8TOW6qbDS3AlEqdrqF8ska6MGi3LK3hyx
DGgo9ocJxBtc+w6R2cP2jWHeMNnscmcee3CNdrvj1aXhKmOjJtiwm4KhsrqrvtP5
52yqDnxFHnR9o5sANJF2AgwhBsBMqBgSctUUYHhhI2WUB+5GFVGr4ETOIaW0p7Bg
Zh8Xu4KdoFGGseLcK7OytYmgLaRTYtlm/kbb8OROaQlF5AXv+lKYjDhfiEyJXDP1
jfH25ardcHFn3tuXY/kr50s9C144gtBPwDe6Fn6AqWG6eZGsuVqOzeaeobbMrO6h
yhbg5lNMkzBsCbrODBsy2YjH5iBegsFrt3aBB+gHrB9I0R6MY97puVN43nxm70ac
yoejTxQxFwc/KFmE0ULtUOdqBHMvK0PoVozPqwTdqTEItNj+r3S5QgB0stFAy3QI
+l65hrZy4N0YMwU6VhM4DDGRzAil8BwB1XWt8PfR5b/ZCRw9aS44xumYW690d+5Y
wyYLDitfXWwYD47QjH2v608ITDF++z8a2Sw8/jGCZHYxVv4MEbHPXD8ngupL63YC
dVVvgrrh6ISagTzV9/GeV8WG3iRBDYfu9kBd6FGVnKwG/cIfvYd2KL1NZHW0jai1
kEZ1czYA9FEvLCmoAcmqS92llFiMjWW20NB6aW2bPuFDX5jORM+j6ISX8sBSy+xP
tAJiy4N5LTwwn2BI1UrRnGaKe9PrAY0QH9uUy40uF8DPno4tP8cCX0l2HNRdbPnH
6G78HbdaP+q2PGhGWrjX/Bhv7/38c+bf5ZDO875sDt3vweiXdzlwu2MAv9ujA+k1
Uz+nkcYUMiHiopKFQaEX16LMfv+h7PK4KsKnhjhsrQjSIuyxa3YtkNhoZ/innBg6
FtmwSq1gjJiCv7o+Ta9FakedEq2X4HK9/FGwYajjdTvWJN3lodnCunQjycL99JYR
Wc8JZliPfAd6VvIttaxKox47uO6jPGi7Bl9dH4OxwFgzjDv86gF0c+HOx7RU/xgy
mCBMwxfuAj8mDDGjSCORNhudw5n39CKk8lvbkspMBWXcc080nOyYquxCoMxN+ims
Nj9ZX1qHxi+0YndKP+ur/gyPD3zu5KZjh8QwzGkoiZdQ/Xerd1KEHNrdhAgLPs5d
/KfB33sxHb3ts+KunM0kEE3/0YWvQRzn6B8LpU1CUM8H+rBVUMsjpsHKHbRQd0z6
cSm6ce3Jo+aFZffD2gs72DTK7vvf8K/d+CmiMLmRNe3GPK/IZsq2p8qVIFTqY9R/
PTStX3Y/OKhdYvL+k0EjYtJgABuLsvXDFr8GzYJsLZ/AxWLR79pdBAHo9CiR8LUc
7tFBqmZhJ4joM2sBW1jCyTgaA91fRBjLMLalvlqeQ7wwdwVwDaSfy0DOQDYD1qs5
T42MdlM0sZx7fX17t/hjHzrkXT+WQMi9xjkjBvWqSo3cCoPZydHGLB+dZUnOGyEh
/U6O2Tg8VSNvoRuZ1pVdRK0JqW8G0eJqMkd4L7FSW6ixE3QXeUlFJZ7yTn4e47Ez
wNkSgmAfhIXToa6JnMXBpsY5V25k2mG7awYUeBNukBbHLBgzM8l4qMWlkQEgHoEw
TLSq3Th3zk4Xv8Ey3UvNhzbaglqoc8+hA+5T7O+kP+3HuG7psWnFVkPSG3dy68do
im19sz6gRbrvZOP4prLm8JEpp/dp8j6nHR9JFBxoO59ZzIUOHbdJwAdROjyw9MwG
rVdU1qu8jZxNRUclGmBIdOgUdt1n5tG+dskwzo3CELqBXcWqCCxK2nS6A/KWNvP2
GQ9RjfFw+yf1WMopamYqZITnJ/4kjo9FPxzhIL8FJk85oRx5IUQjeC2GBaw+gnqQ
iQ1A2SVUeRKoL+Xy7z7JXEP5xzFuUkeoqNjprCt2MtNd/rRW7aKFWdVQb5JN9Nzk
y06xVG+wMADrGyGi1mQYWIPyaaKoVt+JHZNOxl8z4FOKpkPkAObbEaGYQxqN2FY5
INThc0fOrj1vpaj3C23OtTjrhI0mUhoVaTFfFs3oWWbrIFYFmXnXLY+RxxlGWxPV
fEysCcqr5nqIoNaK93LRBH8oSFc/dTXXjzJJb4LfOCnJuCUMOzEKNGYis7MByKz8
UaIgB2O6o28zxucRamavk2eUnCBdfTTj36txQ4qwSaVJPAn6vsTFffPANxN5dmsi
/R/u1hAn00+c+BA4yYr1zABiukxv7UPk2Z8j4/6mgBVjo/HZHpCEN1xzA7pNdwm4
Pgvlzn99ES9pGnoAufin4gXNpeFblYj/LyUYeX9Pbj/xNh5OoN42GOr1BJlpsrCn
AuTvgtGbiIP8ttAKBz/i9QumnyNei9XFy+9IPq0Kh6jUUwJFzJtRM5JxUi9WmqTD
ACisadxhz2KHH+fDCYzHe0dbH8K5MNpWIguJ0mMQDq1tzfJX3a0v7AqZ02fKYFAh
sLvfFpWvb8ylaA/AH6Ysfw4wn35W0dbRt9Hctu1fp3oEebiHyUZMOtLy3DTlgWZf
YhjldFxrLa3PrzOFjFcWHlhW6Q1STUwcJKsTyhv9p36YYY4ErwnRqDn+6abI9h5m
vUtMKzjbL6txPTRHnyLDXW9C/tteSIg71H7ccXuzf7G2Drv0d6vYaKec/HUOZbx8
VCeIa8FtvO3kT+cda1TT03s/VgsmmzFmEpwOvLo8FJt65T/NkgK8SNAPobS7vIWU
FuniGmvNkUbwwFLoupKzkzqt32V4C8ZJ2uTYjlz6hitHXBjBkK+wZelUWgD12zW9
zlcJtkqrzyIoGYdDYAqSPsl5u7IvNYonpRPCPuMCWNtERxLxcg+Ytx5as+H6talC
W3w7plbcS7Uopp299AM10CgLOzaGPWQonpHb5odGvpKlHiSeYgGRfkXWS+OIkPi0
2+rUzPoHQaqBr/BQbKsinywcZPHYSHhNaMkJeGukXbsUnvKGDc3+5rE5c3c1GKgo
ZlgtrbjFZGotlFIdaW28ubzYj917BqVBhlxrrf6g07+vn2tuj3cH9rZ+Ly/16TlG
w/MVZKkZzyQvldIYrxPA0boom/gvwXqbtvxcsHFplZKhl38+ovlupD+ss+xLjl+C
18Dl7F2IHxtUnZhcZ4PwkcBbpSunXmbDF6Jd6/5+cWwDZ9xfV4Y0g8RSWpNlpt6b
wsEuM/bFrtmEX0PossxwL70S2SR2a7YHI4AbMNLBb6iPEWmpH/ieAzQX/jBg+3vV
JtpWeesNUpBseDBEsMNpDhJXL9eV6y5STkBvMTDj8c+IPfa/dTf72Acp7QyEcPgo
ROnjk8XtnUwrNXNy8OogKo0Ix6A15F/W5a+dg1avYBQjd880diUaHwlD0oeW7Kkd
fBwPKar9icswYf1g4UPkACKCIJxEqKZKTmk48FoZedrzHfOEvBD8ZOJmffhR0Mu8
H/cTjKmqO7lpDFhq4eggXHx4BrctPdz4jAmwDLZ83XwY4iRbQDPjNslMwSnERqqq
UQYQMtSjaCAmZnRGEMpzVWqggDTlXrT1zBUBVTDfbCp6d6ip0JNZXBJ1ocNyqq0f
A93V+8uxG7NBT1u8r7hHFnxO/MmJ0h22fJfux0kKxO4puV5t4nsKLBW34wJwBw34
p3Xg5XXuZ7lq7AOcTPkNtYfbzyAU+CzbG/WIeovmxN6NXLmsPzlW4qrjbJmGM8AT
CVSjZ68z668XklCBi6xcInuFJ+wqVXPNB8w9e664Myy6hG9WCjVDieVOuNULY29F
qb1nPSKplEySPa3MVWCkbkSDheeSlrb0ZVITHkpnsss9ha4uj6JN9d3QNsl+aCVx
Eh1A2YTNcW7GeThDdq3PSdwH6e3cYh58tHdPQPUnbPTjKWxkgxFBc4oc6wH6Egnt
p40/6LBAwDFL1Uu7cbUjgK+DenMBE4J1lQjYfMr7prVlkg0NfkvJkAjyhNN0NURG
hcjenwzxQtakRBtAnF7UwFPSHiHokntr3ha7kvYrrSL0igAJapUsuHGOmhkP5pP1
4XTG1bMDokPGBYp4+W93J8qbV9BEhJzj+o22kxKTvHtY0xscOoSw5TmWdT92oLqZ
Dexs+ikPXxtxCVrdQW0Kq0Ez/vZeCQI6TI3QBAlqi9BU2hghjXVkAt4BmPDuYubH
eMtLKwkqmC1jLSm709yAka1rN2yV+6IHjdZHwblUXmickaQCBPi8jYKuX8mrXXcW
lhEz60LoUtko5ArTnR8NQt1xCugzR2lTZdiYW+kudfQ9l4bvAJ3hHibr91rUOIs3
u2Ihp488qmbBOduP7z1vt6YglF8YvJkjMDypD7/TCQS2eSqigyvrmCdwxS/hu2WX
k7Hcgq1S31CrWGgx3ueYxHocxQL6FeE124+P2ajeEft7d3zpfu80lf4NbhNeP6H/
ggFNBPXM4zyI2GeyssrJRB8KnGifeO0EJpRfvxMfGxFemWv2ApPfIweNPO2MuqZC
jh3s/cmE1d5nT/pw6V6yVrd3u9mK4EXPJ12bUrm7rur7yOAhMgbelYaYSV0XNVdw
2Ogn/DBLoGj/GLZIgGoObxMN5c/oOVuYj7Gg/GSgeaVACDfhBjalOhPjzNa4xc6Q
AO6BWvEu0w48asOYbIxW/AwI3fq1IpbsMSwNj/IFnR19zqAz8COILT9wRpkjDMjF
kkMObjiNMetfORfTxBXXzT/NMR5WRK+byvWA33ZBHA/+1/FsdA7FVlUULFL7TdQH
dFPYMu7Pm65j8eZPsi7+9sFosBQkOtEpUTIHG1h1GqeW2EUEFLHnnN12+PKppwac
HSr+hUgYZOZshIjTAHuTyFxc9x7DhSyQ67RjVru0pqmiWOyY3ME0rbmluYo29xIp
0soouLqvPPqJqQ9m5gh/VOxWCdvVWEt33RiragZoZSJti5RKh1JnI0n7i/Xl6Pgo
MA5NRWB6rGpIz+dciHh1kU0Q4nWbwwJj7WPL2tx1Y/jz+s9LbyKQ+c9X+EHj7RoO
1i71lndm9TLuyx6SB4QU16b68DGo9cY7UtJ4vnsGMvgFCq942orktz7A++Jk29tO
ZxFdzYzAVTI6lSReZRQFXzzu1ePpX2VSEb/jyEjhKmDrZ8AId+IJeWuWp0K9T0+n
7BqAXMiP/l4R33QZVrqpw4yVUNJJu+tkvpy6MOZraayRhrj1NMYwJ15tING6CabZ
efXk9eBBlUzQ+cju1x1tPmAWG0J/vkzMuMhYvN7VCEy74/zgabLUgxgKNC60Wik6
Ua/gdMU6ID2FyYq6Z/NbZReNESpD393pxXnMflZaz1TWcxKeYSsG2Fcgqmy8ZHq2
1cGxfWvLaPjGD8RTTd8n7xy0vzZaXwnN6P8brmUfVlf4jl14+l3+s1amFBhh1y43
0sbFAz5xYWfWFnguYLHVwsyIA8UL1mIUrrFCBUG2SSQsfVZCkqeGTY8Sb1Tx+sAW
oqeZmHHUxStCxtbM5APsHq4xDtf1ligwz9kSF8I3XmrMg3IBg5waidgcdo2iwH76
FMAm8OZhBVm1+Oxea2iSEz6dnTn0gVr4DJOYdNLWoVNoB71bB8eL6BJHwO7FzzCo
f8UB13p3fadK8PcCsBT+2Jg4VJAqHAza2nQx8mvJE8XkkbTtOKK/btoAlC+z926q
hSgoyzhuESZbGZ+Bjh4dl+NAAeqeDisCqI4Lo/k8E69mWQ2qnWui55h6F5NI+pm9
5j3K/ZvtOfsJJj79gSJL3g==
`protect END_PROTECTED
