`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cgFPiqhSf+/fU7LVUXkiyQ1B32pvGpznd8Wuhd2mt5Z+ZiCKIqXI8HZTPdRqX6hW
s/lz4cKbaWiSpQE2ylKpPqlA/YOL55CDgI94jFssJYRPMMn0jg3YeBmcvpR5DvFf
fR5aG9SFE0C/13ohceP4HD6TOb5s7do2KmkW7PNDR831vl5Ls08ebk6boL5oEoJx
ZpcSffrNVyAH0PTQZtTUl6RKEoXOUw9DzLCGfwR8fddEGz2w8DchwpJfbGDCq2X1
GZZM0ptsSGXe6Bilqp8dNFGipwjJqE6RWAC6w4fYBR3weVy15p9behX/tLU24NJM
ZTnmUNvtItr8UfFA8R4xl3KpQwj8ZiCaIXVl3I4Q4K7x1k+e6PD+s955WF9Fn62/
opepti4TVar52XzO00p9IYmTe+QpjP35iAhklUz+g0+eOClPdnSKGSQKayYQ/3Ua
jQbqCGZStztd6SgZNNKC9Q==
`protect END_PROTECTED
