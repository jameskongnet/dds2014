`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K16CGA1QOSIfvgc9S1wIUMp+XC6++30VLBYlOUXZvyYIICtRLtaxzzJ/FS8rwbCI
pOLYL0RPBINLK+fSJtnUqeHjqDY/fllbEESbtbpoKy9rVtWab4+qaWYYpQs5Qpmj
xEzFFDI6D0ZsSaH9dIZyTl8KL4L5ljBGmIxzzw0eTEWphXc7/CHKiKALKBX4FqFK
Q0qhlyHe6waw+GkqlUONOCbN1Ds6iCRn1LlLyJAGqT9nbewjqLTvy6Oh76u7SlzZ
sbWul3PuMnA5Q7PKIh+hbbLoku1ej7/X+SIDStLNRFahwiTs5+m3KELgIwl2CbMQ
Kb3k8RR/aZoim+vUaFgFyqWYYUS70NGVzDLsHgLHHvVR0gQnnso3bSDfut2JEF+4
hKXGYakbD62PCwbZdpaE3wMZEUxQh0cnEZJA3XYuB5fnPf3jG+0Z7A2L2DvuxaK5
sTseVWEjpYVr7RzOO+O9aLQ+S1lFsB26pKAGm7phcy5yifUOYnTMVaRDwNpNdXy+
e78tqJpZZW8wAq+obN8IZWatE9TxRcGXPnnJa809mblgVyyK9fiDxTEunC660eh0
fyHmATvRt2nJ919lvkWI5QPjbZ/k1JnzbTws8UfHo41K+EnYNIDxknDM8vpvki9O
GmGLx5YSrDRcfLMQ4DyRH5P/tuJzmHhSb4gz7eCLSmKmL2xI1HF8teES8g0OcnCk
q6gNiqL8aQE09fGymiezwrzzhE6dTjKwBDs7qiujFbzitww34i7wklV0kQYM2Vux
W438aYTzygD4zLRqa2m8oczlB3WxCqmqdhGzp/cQZXaufvpxzl8eGKjwrWng/khp
AhFNSmDhuE+ULNx2vcHEno5Fud8gVMq80cfu89/j6wnqUg7/eA58ECbhyMBFgjNI
QmiDt6zodBbnd0Q2Ayb6uI6SAw63D1XaWphZR21Gt+8mtdqdu4kFW5m/AhYHgDb0
SqQnu/pCzybbU7V+nR9xs1WOV3eKlLn+x8uErsnQMXmPxy4amwl7or/FVyzpxtPR
YRpZnHd8vMaT67WI0H+swajm6Gl/rypSAiYSixxC2HTKK1kg/9mA78akSaGifsOh
yCful69E6MsDx1nqtnWjwLoFnJOoUnzOQDT64MTkkcb0rdvKaSlOBU8fWPBx7chy
XNVpaZXqsLe1BIZntFu6ySA1aLkKvzkeivE66PBLDZ7YkT8N05jFZyIa/hyT/AvT
2/6CtZlXUdfhZWr5Dwnjfqn4m6lyw8fTc0EWjDiWphDCdq0M69HcwbMD9DN/gmqr
TDfXOHSH0+UEycHBrXF2pWywX60lRVenZK4hKZ3tIKPk4Lx9Z43yEKuqljN87rm3
iSrqlzIotQx8SA6nrfKCPfNUJ4oYGw1D3+9xIoDpY4Sr+Lbpzg/nl7UJ0I2uOX52
QsrQsCZp/HaHBgl4fNGzM9VEj8FH+2Qr9khbOhfj3VuOPFrsRYo9uiSpi+rmIIxb
//vEslO+4wfjIR4b0QcGhoNSUc8TSq9RnTLT3NlNc0dDGINfq662fJoXt+qUkHes
oSPZYivb2S86TdUVw4Bky7ODu9DYp6HbaF6/Y9uFn0tX/PgHkqNv/aMF9jsEvexz
Ov8lu0zy/SrLs7wt0VXzafe2rWiQ3Oz+08mGTR3nDmqA9OcYu/YfIemEPbSPmxM0
S+vPr6XHYavbsUgTyLAzspOuG1FCdYjoFeb72AQIya5a6yK4sumy6Q3rprBo9pwz
zeJFJmMcCR1tZogAXp7l1J6/3jAX6tV6bzen3XFapzkud9bEk12GQWt+3TNb7k03
DdbV7IGeZzm97XmYxhY41FmpGKiQXIW3A0gJY1Rf6y9zZjAIkNp7r01eX65F9FWx
j6qfd+d+U+JRZ7gbGgtE4ydhpnkO9AaLnpLO9tFj4l+2FOwWPJFKcyh9z+qbeiPQ
zr/a5TxYAL5AoHKHCn1oBtfCguqq3OPHI/B/lCG1QUjFJ4uzmi3nB+utGfv+2l+O
6UCXQY0QbY4uPbqO43d++m3rV3YFcWkpiHAKODEAA6aODh9+65hvnup0CDkDGxeZ
zZ2uDAICD8EbvZpTOeO/Q3x7HkrwTqXfDaHDsJoQ4u1Bf7LMIiWG/FL2jmL5qPk1
4aBVZr3yWqwnNJZF/UySvBnsJNC9sWu4C2PnOw1zg6r6LX1olPwl1zOeIThV0DUG
eSSpdUZsYhoE0gaV68JTVxlYtJyH/SfcsGOpElmryK1Xp19B8+OU24FpctFxyAe2
fGlMmWX3l0oT1aBcbcFTu+UMQrWIuuYAI/kQnJ8MpkFuChlaiULctrY6z8AAQtPX
E20M2F/1Hr0A/P8amYyVIPIIyvHfWdCCwudKQo47Qa4kyPpHw/lDx82ivu0XkB4c
RCF3ANb4a2pNWLz2uCWiH1xXYwpba4TgtoadnoTTQqfbwAdPGzgJzAH0YO2/v2WZ
4nY3dBRu34kCg2TJ5ZniG8I2WZLM5gLMjaKeFbwzCft0AFkvNrWq3MF24naOJ68i
Y4HMlnt0XvHt155thIeejTgwGFKSJz1swhca3kiULE9rv5/l8HhPijjUGKh8CXm9
uKvqZZeL94nGpTE/5Es+bcIEPT0QdVKc5J1+36jegpB6xuovQjeoDrXXvRvV9UzV
pIwKnLsb2oSkXntGK9tGyrvtXKa64rxU9tMkdI83HPwZTiZrBj+ITxTiMQLtqSMq
mpTmHBzd3XnrUubicEuvkrV0lWnUVRRRhpbb6y2XqHeX7mH7tUivy4O4awRJDAR0
otPfJLKOOkVfvbOZu/ke3gNXQSnIHa56lvxtrbLhZ7Yx+rvmPu4dl8ucL5Pyv46F
7ogtnMsMgXFr94bj4QPA23glppX/WLVjFlboHkfrcGqrl7qi7tiV8gFsO//00gHV
b//DqILtjBq6M4B90M7TWCXpxQ9zNEI2uc0FaTd6Gb5TXUMoeRTC+3s0DF35utdI
Ic44MxtxAEeUil86hRVMw9WyBRM8inf+wXO3ksfD2uYOpKpp5nbwMKstr4OtbJZx
zfNb1cPHpdhLHoLeEnSw0vZIqpCQpNxC2xrZOOYlJTnVXTVexDKESWTUuaQorQkZ
H/0eAsoqlICvpmpvKvASxcpvTYc/UX6FC9iK3bZPtj+Kkhv5862vkw9IBIaA9dyV
URUWlk3ttwM6Msi0WTrlVo4vxxLfRaInZBjIHBifRu5aluNdXg+zx6uDGdXnO/f4
Es+QzQT7egBpj8bdz3LlEIz8cYAIh4JEho/UK9mkGCeY9e5g+ymx6qA1SFcS6AD3
KePDBAPiLFhRxo93xssN6x3RCstnv1JrLCMJHr1S34+m0BjZSC/QzRV8j6tL1sLS
zg/Z76uuIQqNOdbpkDzfj85tu5r1Gfx8HSwRRNx1WXHnCoaEMwp1BvnS/5rk2e5V
DsL9xSHHzwFVeqbg81qR/d8eA0moALSc/rzUskIb+VubPzC21YtIwsaoyga0N84A
kHJ9WvLLaBRK577131FU1klAmr05R4stOgaoPC0QEqa79YUO5p0oekIZoh4kfYwZ
s6Mfe16QAgerNsXeu6snau4RTVeqgg1dlOE/BCNVHAUwiOweNIV8olLBKGwISG2f
u34mlx+7XbrmnM6FprruJzrb2kp2lRx8EwNtrUFLBIyc6rN44oNpIQ4RD088EfXD
T+qJ/PxGK16Dvtuh/L3ty4rzfGO4ugRoeVgy1Sz142dvW3SQm5obvyQ8SxDb3BMI
/Z/YOb4R4YhznDmP+dSDz/o116sseEmYk+/Rn/R8iTg1GyoTTWxqJMSXlcfJKthj
2BT3BfSrDwden1pkBbghLFRSUGU4MsS76NeKwUTvrm5KvdY5RXKQRL0UIxnxq+O7
RbTYKjfikr7yf+ivD8ZcS5F7HnN3KlboX/hQTT/wxBvA5GLuJY+YGX2zCi09AiW+
yza7dZwjbYmqhOPv4+MdU/ZW9Vc7clDnebbKEVFo2fHuEk0KLv58Dr3kVJzLPrpI
+4//o7WIYRkmBc+Y1w314D3erdjIsihJ0Ol5U/pxSSGmPVPT/51wPg/3fAc+D8Z5
0jrQXOE4MCZmY8AKGSrkZi4fdgxcbrMQaI9QxmX7RH/7j24uZwt7Eyr6Pzuz2Rzv
VOWnvyh6SxzTyohoxQ7/M69KJetWtpkLLd7BT3gQXLnxOwtIAQKs77mWu7+XaUN8
mwupl6saSzJQt4r1YKaDm40UQc/2hQyaMygP1JcemUGX9j+2ra6OyLXXqegVAaLv
3kFCYvbFYbjqukHeZ6sUyRYbGD4c9f/y7YA2w9WfSyRE62WWMYhiFimFRZJXGk0W
6JbkafjQtJz9xwME1Zq0LIJSy8nbithl3i6zJ8HFRvH67cC8A9NxfAHEjultjcmM
MCVN5WjImuACvqzJ6cuUm1ILEJ73AYqRTDL6srWpUMw17vQuFsizoSzU82CYBuC7
n4rzn1sOk9NaIVjghrpkt3W+bclAKTPeMge7NQg8Z3svsF+qtgKWRAeGasDPAub7
AhgbW4mAgNrw5HJ1otRk2nJfx+rtuQzcXL9FNoxe9wSra4Wp29dMLW98T+/BOOPf
vjgXEc2TEmu7FjQ07Df5ZWPeLrQfjsC85fEW4q3o/f56+pF0fjNeoTI6ZnrLLV1L
xVWBY0g0iuzfJdkNPCIezjR2n8R3AcqFEsHNozxy228H4V3P7NG5S5FeUyfiTe60
SXc01iDNXAlec/rEZJ0BU8DvHiBZB+Wdk55ltpHC3QLNZuccKP6uIA+MZBTLvnyZ
stwVf6ibtvTugw0fB+hCP88PQnqOCsY3LcOHwrclbn3NGmgBtrDVRyWywz6JmkjE
ZzDEC0EfLc2cyI1erJcZ5Ny39bFkjzAJmSN6aHNKZ5CgGDhErM6rSQAeemYfdxgV
uL/m4w+ufB5ODY9rjkoXAv5P660AdTmi2f+n/PaC+MP8kwg0gTOgw3EDgDJ8YKKF
RMPQUn4cpi7jXG4rZ5q8UuC83GrCekbWcNkJGyHSBFlpJ3BgF24GI94dFkFWPNyu
BUnhKttoTyCwFQMtsor5R0C3iFlsztyLluecYOZx+AmmGMM843aRtiwpWvYkXR3y
oWNOysj67/XOHMgQZaVEGvEb6uOjqC+tQfq4s5Fq5tMevss6ljQPfS8zDOdNHc2f
Sesymeox+5cAxmnWQd+s9Pr38wdE1/lHEB17Ho+1cjFLmSA1YKr8PcCAh+MwvGeJ
AugnI4XDkj51c6cF9ryFaw3Vklnm1PCC7k96v5CnPJFr2D4CX6FhDo2Y5CXe/+kk
L366QcumUS+KD2npJeH7vgbGUAwfxq+TU76zcNlQINpXx53BGc9Oe9FBnNoj6bOw
2BYQrZozcprvirPJ/flbZTiyTqU77LF8GgQhJlmBdegmgyXWJs/sbnVGdgdBsljW
owI/D/oyY0A6tZg1Kej7czFjhhwJDbTFYOG4y3QGB6VY+pzG3heZJ3NX8eNI6CkH
DOyThyUpClpsoEim4KAX+rzkEz7ilkyJf3mYJ7RWQoceFnaiX10yis8sajXl/Djj
+ppTTbcHiJ5my9vSDFPXTj3Q9pNuf08xyT8+lA8GnbkhqCx1Q/Q20xJkOS3ZEwtK
EV0wB4T0aZH+KeNnaFI6FL/uwB5eoBxv5imWLlXDwbQhdytwNE3dksIz+Xek0P3f
IHeRwwuzhlSlsYFhxZRacpUL7+ApP5TxJB7edrT7lwLDKS37+8s1D5hbQ8XcSvtG
+vp2HQwLscuZLj6m3zPB0g2Izh+cprtiTsI+uxp25YJCMNZfLcpu13ifvwsW7mwe
sZFvZ7KE8OuaLVrUlrUT8w+fQV21SSBM0Lm2siqSZqpt43OopcPeW8kZmDRhPv+m
p5a9kulH8K0gVRrSWTZR6fr8XKBs+ihnJeyU3TIe4pe9CMiCZL3xnRpB4W12wp9E
z8mkkaf0ycbKCI+pXTJM50r/ArC6Xn7mE/Sz6DRkD8YWTF9gAKPBhbBiTkXumjao
45HTh98cp3paHqZaHFpH8MMdC/ggWB/kmZrGkdXeBcXDR/HAscaBYox1eeUMXGdE
acIju4nn899dmLP49JuBAXRtWNjkxvSFcrV1G2/ogotdX9UvfNbFdSVm+naeoR4C
mjGQ4VFe4s3rsqHtg3F+IWy1/FjqJMgaivhYrPjghw9mL4xu1aI6mCd04A1vBGfB
D2+518IMD8f0zgfYZ8UBXQcec3IuUNSxRaXj2SoZYNBUiuH2Q0u4aZfwyp09xwds
0y7S/HIg0KveNcrMb76quVvlbB2HvCnfPhGIjhuWUedrwderrrjM5h5iR+IjEqPW
004zn1AZKbt5CbVlA9aRTvtCWKDAD6hFjBU4ItsgJ62TDYoA1Jik4AOzD+R8rsg5
UL5T/jaLyPgvUrRqSSvywfSGAe8i5O3lMJxmr2s6TcsRvswpsekblJnc9xFYXrzJ
z6XrtZLbBFZ+RQDTmwmLu01iU4ILe6ZuNqzhUO1Ozft0Erx7hLCTcAxNSg5e56NO
Vvj5xpNRcsiuUCo2JezTlc2qrKC/HIuryRuHRXmjYcaQy0NCpChVOt3p8b4747lL
JOioyGh2SgLqhmjC/QnHFSMbUkN+2IXInwNd0tE5EJgM/IRLB8hGoJS3z9pK+pOW
0lub7Aatov3E6upOnEUNDqjUo5LhuQnVC7a25Oq+5v9iOrEJ+t6AMSTCUQUdn/Md
dePyDv86poeODGZklnxFwLR+hLs5zm0MGrD7CHEmcT7r9kjc6skLvParUIrYxRRd
YTZYSn8GgWJQjqorFMAI4Y5wTHwfNaS2wMgkC02q9HzWVceatC9LDHj1uTHS+0RA
ihdfa0C1CashiFsLMo88jjiEAjq6+Zg2B6CowYWyU4jwN1l2cjUBbnUOEmbGMJUn
+cEW/XzTtpzCWY2p0v61+oQh9g40lHbvBhsTXkhlUM6AU611UPHX7FOQ96sZZ7Kx
8TERqfpx0VRfo41xXiyqYRarutciYzAf1sdP7sLO7rwJSr7EXKgant/Fvf9MgFFx
MlIRgaVgIKBP+xEnpt8QjannGuKirZhnPy71ekbTkp2vDQr+p5/aekwWLnLQWDm+
/J/+BHI2yqpXq+50/SsgwyxGjIFS7YeMq04fHg/UIBcCUv6GY2zk8pglXSOjOcTL
9NMNYLr5btIj228qUJD7P44eocC4GTh2wTJSEMrjndCaU4ca61y/fEm8vDm25u8/
hUOSrrZxJmN0JGZckPLqFH7pzhPM1lZiolHgAjnM40VNzF84KAaLpFOSnyT16XVf
irQGAEvX+qGyZU0aj8s+IrfPvRdVkkE0amA3t/nPZj5eqSIHJvrh7yfASPqglGI7
CIzM+yZsvjDkqj13oSDW4gfw6ePgPdxcv0fPS5N1rtOamJ3C2WRZSBSrysgffA2T
scinXihcXcIRThjLseqYypcVSR88SKDeCkYld9qlLYhPJRq1Er4stXcXAELEzquT
jQhtkqN8Ku3veB5OD/87jE+bBIQtDtg5zYhLTeZXN9K7dq0g/+1Ns5vAMX31m52B
TM33JEh8AK+DvpKSPowBXg4QBwPQsfmpdRER19LJlI1Pr75/mfxwY3iTnJ2c1eT+
BlOXG0L7XKtAtBhS/Xa7JvZ00vLYdWWnqOFx0Q+VDhTC4XcVn+n9kYMJkB6MSyxx
Ad8CaC3vgVe7xrez1AR7+UXDBNqC2mj1hTZOPppC/GRSUidWz5kxoiVrcWNnmfUa
Oq7+/H6WvkSdkDW8PVQwp1uyj+63T3AH3+h76uiXRuODacSXMYgboIr0yl0ehPk3
aFTptIRCCRLK2KzehcCyKKIPOZk0Wl75YPyFH8PwBsn86XNAy7X2mWRVD2epGO1D
z+BAxM/DHvJ7OIeL1+WFTsF7YKlQwJoXie1DntKv+GPfKFC9ocs4kwFtbLQVtJLP
lQlssZXYWGx+QRanC7bRAdPQlpOATsdATHvq5CG1ZGVFExCX8rrWnAsVsXK4V1hH
MJ6aFMqHd8zPDeAYPs4s124Ms3yUZggZPhExOhdSnmZaixe4UjjNQhRajI6VuGii
bHXO6g+cD5WUsP4nE6vBKbs6HLH4J6RoxiKWCwUj7MJ24ihgFHCi21v6rG8Iuh4t
TYCSmtPQAnAlfUIGmh59UK8i8QKs2g8sFEi/NeUkHdDPfR7DQHR5uxY9Ve7ZAGty
hlKyoD18x3xrdNyD0gl1cxYh2DmUNPUXtNI9exVqH4pObdwFrAQ13ZTZGFV7Wd1C
+pl1Jy3cxzjFTJxqx0apx/GJuaJMJBX0TKbyAQe4viTZqVVQon2IAhao9X6bQLtg
v31NQ3bsmkGRQ5nCrKd/tSyYaacPXp0qRQxfvQEnGSK5HLbuLSdq6QXQa5UASJYH
e4R0E1Yu9GxSsxH2ip2wDXsd2eHbyN/3QdKxtjmlfoZPWzvB1Nh53fNmQ23KdiZj
Bj7mLcmnQzCBY24k2lZCh/DIb/QS9Dmmfw7L8xc+YH2lwbEji7QCxMq5o7hK/iaP
qmVyRWT2dCaXK5gYor2iuyPscCs82EzF8Nog44Tf/BBInIzXh5yVMYl1I2GMJJtM
HdX1nBSCLNPwpTFVr+RBqvV/TVJuwXNoPrnsiyBS9xOqiOeNZgkwbCAXw5a27vs7
A+NVynU5wgMLyPny2nECXcPm9kpx6vBAXUx1R3Cm+Y1xaXoQQ8KWDSws3qiLgfK2
V1YmLl6rl4RlDd0Wd7SF7PHhY8acJ3UIERs8QunkbBZXgdfbB637Px4R0VGPl8/W
Fjz3VKRhzglFce17r/oMwGA8dpXNb4W2y2MIWlPbnu/rHDU3Xs+NUxq6Ct/z4geN
cd9w56G6MtjdlIoXY7bMLz9XVVAPDPOy7LDsRFKSW0r6jD2XcPlWU3lOu/OYaYPl
xRmxmNYKygMr8vR7HK5333roKoji5oTiVs6KesW7d2fZ45Rf92dZnMeOWgB3yrBJ
KBQ6cyU/BGKT+DTsqHeQkKBekGyxm2AuCTVg6msV3q25IBMguiN8j3n8yhY3dmjx
0Hq2FjW6Ggd9GQb9ytiWS/G4paaPew32ANIdnwV/BiznZqJ7x7IOMlyXq+rDfsbc
C5uldwwh8PPMCGxk/JSuChmKoeq55bvBC9lyGpLiun/QiZZJfCpodr9FCFy3Yw+O
BLdpUakSwSIGAVvm0zSMtRYxqrownwgTyIz5xpDeGZ5uQ4VY+g83RvlR+VEGoWxc
GSwD9clx3NLGNU3GzeIaFqpyCHsbOXcqtjS7mlCpT8MU+wma24FOGc5wm+oT1HRI
PSBA7yX3MH5CwaKLc1Sc9NBnLQfmIamOayJVjDoxxHE7vYTJSXetks6Dz+kYzoa4
rx6mBF7z6PBdb57vCQ4YrDlxB0LFmERTOTrNS/2py+kRIf/WB8QdCfVYhi1T42D8
213nrnJya71Yt7XohmmuP/A6KKFiAesfXk54WoEyx5y4ddoLm8MpwTt2o6QLh842
3oTP0NQONnZW2yXb3Mm+W8cYUxB9x0yYl/XaAmnkp4dWEDXTHFfRSuUvZQb8yq1n
ZF0JNTX7suy+NXAauLXygcdCnl9d4n6dO+WC7J5fLSwc/8S03+jqlyJCc/IP/XZs
o9Crx8EsydAOOTneKYiyGxdGi6QtECpMxJ95WeCKSLL51CV1GATtto1voM5vWLSM
OFit0XGt8TJ7ERORkVYELQvpZEuC6LbGUFms4oG0D9x3S+yerRAwdJf7FY6bUmhl
eXijJW/iPOGYGT60Elhi0KDuXgsAWvPT9YS/6FXIRTYBXWyrvqhZq05aReOxzEWY
c8oHemotz442Sfy6lNXfJhKNJc6rQNUUag5rDGZ3r1h4iMPg3J+VM6riS7vDv+WN
eUXGZrYA+dRX6qRp++1jfbW/VZIZJSTbB8+EyuiA/ihTS15lScFHoQegqg0W9RxM
v2NOmzjGImvZzPgoRgohTQ==
`protect END_PROTECTED
