`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QVnyvfovuQyPfCb9dr0OVkI9UiaZPb7PdjJ5bTNs3bBk1ZLKYKG8ICX0sIZ92OyH
ktjJ8iFtUITux9U4GHqnAwmFPR1HVVmSKO05MlfE8p97CHmYhaAr5Vzj2fWIbwSx
9fO8qwdFWWNLLhxnLOODnOXY5xrN4YPBFh3ISPdyS9Hn+DTcA6VQ98c8w4dQD0Rp
GbgdtBafjgOldfnd2OtsC6YXGdo5fkqY6f+vJWYCx85zh8T3EhXZxXIQ78dOU9Hx
CxA+AJ3u5xoB8fwAdWePmTsaCRGgtPWRJclYxeRD9vgGpQm4wHdnh4MwCSq0JiFq
mmrUzLKi7ClIVPS6GPHeUJ8VCtvN/VtoRAA/aTzE12mdscD8Bc4chFmA1lS5JQs+
XTTUtKso6y6vgtx+3ErJUQVYCGHnDmkf9hBVGA9HpChmwGWrgrpWj/QFyPV2j2OU
g/HYAj7m9r03t/7niH3qRV68tmt4wA08CvlcNeua05yGipFFIAx1JpDLzmK++Rxk
aieQTs30wD0+cAApJ53m8efNq7C/aGtlBH1wGJCPesYSUsOH+WwqbxcfFd+6t9r7
0TCJftkEX5Rd+TI5EzReEtBiG35K52okPlje6X/jwLL4IgxJOPuwa9kLqt+Btvry
YHlSIndUZ+RN2gfHABCuXyo2EY71VpDwiiin1L6iP6q3lF1svwjHuW9Ma8PnNfNq
jW6ReNkx0KQhn+tHo8HQXEGtrZ53L2nqbFcCUAdCr0zwL72dwo2+l/hKOtSWNBRB
+blJP0ZHjra9NrtNGaoZTjw1bPaGtHxzTi5sbEnhnfgi+W/d07sqpmKh3kPLbfys
Y9k2BtJXJZFCcwuaCF7lAG8p3PH1wzupMcezBUQyzH75v0rue3ifMguqm/ThFNKp
HNtOBhn0PMbB5ZfNJm3DJHCzHRKd+TGLRgjoFO4NKPVNsO2MHFxdVbo5ScskeB9v
UGaiu3a2RPSZFqJU6QEL0QNk0Nidfq/j9juhspRUex8CyNogt4hxqKww7fFoDZ7L
vm8SXOnL5uuh3xIeuvYfd8XdVFzXxYt53tTQYIQpEXdTkE6vOO2sEyMZPrgwsSk8
3VpniQ5ZAtlkg2xjlqxnfgIsJwbS4BegEH9tww1kxaqpzA55tt7tazoXOTO0A0li
RRU5o5FzRX1zLyT8OL559c8CdQhevORx+aJVwJv9jeHD91SR3XMLlN6Rb667K+jw
AZuAVsW2PKwDhou+qgwxiOx8/EBCk4jJt/mTo48FwtwkisEqdFJSeOXFgN3adkxe
MYLsqNzvbo5HxnvBc5kxjERP9vmPC6Bu95T6Q0K29JvSNUZzKIuSzQ01I0UYqeF0
SvWurZsHHNrIAgZMuj0kU6ux1quJzSCqT60Ej5lzvcq2er6DN5sBr8TXxUhLiuJ5
WUR3CEECA4e3ISTb6uKt9YThzDH/iI1TJjs4DCorNHOVrGNB3LKW+XIYkLlPvkbT
QExdlGnS/Mrul1L22DNf7eRf5MHVZIxHm7dSNULS8scUStDrmxOFgjsa4Ojq8D19
wCRpf6wWMwEVrKOvzldthiIye8zLph5XM/PfEj93QNGtpnDueNns5dMwehhpFw97
dlhL0SMB1k0zvNja0bKq46Emg/drIKjwoLLVwguRvFjFWqPJB2OyfWaMggLAXMm1
F5SUFvCnV61t/3T+bIqbwp+4Zd+/YoZ0O+3jcn1cSBRVUa08eVxUWlx/YlS9q6qP
eH3QeR5PgztmdJWzkTan8WriCDJuNOyGO0fuq1TEprcbU94d+2JUcIzRr5moa8nr
ngzjNOIj9Fe7n2CfI+RxKkl4jABkqfWXNOmMJKr4ZYK0cELqeOqz/NyF2DU9qtEO
11fQYBwFyV47ott3dXJnn89f3VTaPvubPUqXg+0VSqsPMhxQ+8v6Z41YLyLUuh7k
OGGclc6/5kVLZVWE9l1LRbdZOQy0KXJ2oHvCF+oqz/IFeTbYO7H3zhHHcusiybg2
CXroRPZoOGk1QLrnYODH5oIf2Iyvm+cVS/ubXJDRh8bSQIXNYthPaLuYKGZ4ciQu
QcJf5S6pHRvNfu+xaULS1XQhDSZ5lw4FfKpb7oWfl4345U9qx7EPvQJ7ucNSHGvI
OeJJte3vmLSWuaLWdjXYdQQl31MfNF9XYjlzRBgwu3RF6xZsv13BlqvSvaMNLdGD
sjEVaYPWlpHpshDKKwTkyJCc0WY5auSLREYwHHMsl+TKIsnCW5nHyeKZV0QbC06U
GnkhZMn8q820sWeucvvnDU9B5/3+FhkSRbCYH4iWLUz+KDiUf32zjgyDI/QPd1hO
kbzl/WPtmSrPOmIsrRLC39lFdocl5wgRJSKPtrFwARQ+qZOfoCSODu5uRuxx1YNS
Wixjy8/ATnAqjatGDURa20I6NSnMzMyBhWgmTWSF9lU1KQy6/rWsmKKLqIJJM5lx
viejFdNIfVGPCbV3d1NRIW4rcYSDuLzvEDx4mE5i2urHXgOmj52AOcUDL7I5mseg
laVz6QughKRGPBTbymQN1MYWL4r+LKmz4Zni0RPnzcovrePKgyIKKpqhqiSOS2ll
w0MoDTTeyo1OYg1+2LtlmwLtTYRvkAOUZVnwOq18jJWTz02/Z54fSyIK9MJK4usf
UjZkYPL15F9jGw8aXfrQvn60M3/UwiE7U9dYzHGa8Yj65zOXUTwWjoiOGsbykR4k
zSz9tO0QqmeCI3iMTiLkmsBpGsH+nK8DeySnPnB6bSA1lUhyIScYM+PapPFJqAcZ
a1ZsGa/UPo/lp4Sc0SxOXmMi/ub5adw+qDSACCu0D1zQvOFIcmwXobL7knGQOdMo
IsBuKRX5qOWhIcxxWt/OWG2z8JfGGn3d/5jIXtYmbs/1JFot6h/5K61TdfJRP/X5
E4mxgosElSTRSXvfL6PsL8nVEAORwCL9abaxXjmEbjarM6tMgvIdCAOrEn/0X9N4
CMlBgpFsiWTrXlKoj0B2B0j2SLcd2jDWHoqdX4Zbu/6VDgf5uOwoASEXd4WYOmwa
xKl8OplcQGow/ADeK0s9e2nwMXbIaRe4gfQQcmKRj4I=
`protect END_PROTECTED
