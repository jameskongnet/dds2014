`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P/EvpZtktioLeWgujjSYac36koJ/5itgy6xWmdkQTKIFc0LOT8mZv2l69WtTn8Aw
yqjYsW730jjQFS+SXJTWGjPIxL9ECl+QYKvTMJpZVjKwUTSOWi5Sc6PMkvDOKsMf
wB4xEPKk7tJ/LNIUy+nAVXzMkTuvyFR1zIeWnGPLPcQyizOJI4iGd2wlbEDg4Dje
NRi6Xld8nTX1NhZWpyFku3ktxcgXRyKeqhTjUwsGS7YcqkFbwCV6nFMxBWUejT2b
3vk/BQbd+aXImpTqJm5IZ7pU08BDa0acXraSg4UiphULa0TQjRmeIanC0zk/r74x
mlcz12eJkJ0s7JDJi+XZsVre0g6pGeWxw0Y2oSGHkdLM30BkvRnO51tDAZKenuMh
svws+qCaf4jLNhQkAksUBRauz98DSQZoVI4z9E7fTXvSyndZFWx0N62bfPVoUfNj
yIwiSGJRiBoiIQpMiZX+xF73BaICxYESnanyZ4qaRvTVJzTb9mtdOQJvOGNnXXlX
TQC2LpWcJDnN30rrafEtnf4buCCgGEmf9zhQK+snZ2OCab1aHedY3JOwsC/UHE9I
+d1Uqv0TEDXvjmhRlbA5sX4R3w/y7SeqrOhTWx/96c72piHBzkn9QGHGuvucOxwH
jpM9fI4P9GP0wdr2FPFKAV6vnS1bMRqCN6+vwP8lRMkrOhvkrWt/psq11PIVzpLO
uhnXy9KFN5m0MdyCT3YNkA9WjOAhWEXqm2LYu/vchLp/FQ2GWDE83ko1u3NUQoDL
wreBfWcx+yCF/jkN4mZGUaD2h044x/uyajAsSOpCnbv4R8BVOMyxN2Utph9bBEdz
xgM5fLkqnlDNXPSJ7Z87rw75Ny3i852BKrvAQpE+m/Vw9tYib/SZwYL+B1r9STXF
xTfd5ZEdHaguZ/ujsGTG0zQ2Bg2ov9Meo5FI1w4SB9ScOWeKOHT5cnp3SLBGFWdH
4Yy+S49Nvnqz6cWGnMNNi1uxYwGJi9knVLN2ieWlxheXbC37EV3AKyGg4Yc6qgZj
e1Wh0xFmo5tNPd4wxy0WL7m+3IrAIaKpvJ/iKaaa0gzWszZaQZVWrV1oYqW5UtZ0
vhjT9t+pxKiuZVjx0r3Wgf4Bs3Q8fZfU9d4XS4/jqtTjfIx/VTSWCFn5K8zx5hak
ejRLzuzjTa8CsNOGyPPs92S5azUKzvmhSv8ueezezW4=
`protect END_PROTECTED
