`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDck5nLR15Gi4ziHZDoDgUOXYxDAKN1N/bwW8RGYGM6XPOiJCsah1zNW+Gq/GkPl
b+3pADKYaffZ1yNBtki9eNUydp3NQuf0i6sWea5hf92vm8JYqOJrLgnybtGkxddQ
HgCVu5e/yxnZI3iIpwg3HKaTfeKQWOB+L3CX44WbopNxG9Ff7bSS2K8RVtD1ZBZk
cRoybb65NEmYuY9J8aDzGonfNvCaRGBtUwm8Dvzw5KYW6UwB1PoQk0aFie8VvXwl
lKLaD7UByyLkBqQtOXbEHIpdBkBa5Imhsk5o+pzvJDhGTMbfL+9bJPjrBzX+gjIa
vrkMG5owI1jSvkV1H++LRCnb5/Q27ZihMEv37A5m+NS2dtQdb1NfdXbClPKl/lO2
6m4sELS/tYhqjaaNomwB7eTnXivd5vvxWu2nHvRa0ppQEGp3klqg61WrM7nyGZfz
Hh740C2SLBd+Tt4TwE3MPpz4bkrY7zMqx/uzcTuIcrkXvN/9Qm242HsTVHx9rCtV
GBMRjCAynYSAMZIRzb1mDiwnE4bSlnrbXnXv6k1zQyM8SbIcmhgGaomoIiIqjsjk
G33fb7PEyIeiZWed9AXiRHwaWUWlfBbyxW8nFdVrOxB7pc3QCydrHswQXH/w4KsU
8KB/V7Ew15tY0doEehPggmTaWMcx4Wnd3W41ZZ/P87gXxNhk4ehSaSByOBKIFfqZ
3+vVxhH/cFgkyv4Gt8LjdRWmlYB0rl8ZblMQPoXRiL2QNivNMlzKatzNyt5zgCCP
yu5w347jrDpU1wDIIIb+cj1WbTOq+sk20dJuuLSrgUHSyxmSgBFnm/h/4jveBXkx
oBLk2iFNPqUTN/yYEfqG8TI/bA7IHWlfxB8Pa+SPL+Ub/FiPRBIjhmcHSTSOjFPD
CZgUn/AkqVHMYFt9Ji9kIk+EqSsultNBfHGMkxip6mfrXV2hQeH2lmpRgqYYKQHZ
FRncA/PUSOEoMZAyM6Altu6z4Oe+XuWVJJOUkBvpgh/5FtyjQ/lTJQ0EXiZ2NBlj
0sFmI6cpGz2Ktgb2J8kLFqhMJsKGgUdNGT/F5l0o+agKs5iDFh4kKAGhfSjE3Pxy
Pc4v5JplFXJ8XvUHixvvbcRypQev6LOlKcaa2SawpFBuXbSIL6mzPcmr+isDOiHB
FbjgCEb+NjVig98dYA53nHJ1IRkAlINTqs9d7Zsmd5p2jlffLUnFRuhiAg/aTIJp
OQxe2n4yjbxuyM2YnQSxQOX44W/vxQOq8y2ECVq+UVndQC+vXOfJVmx9+J+hsedW
apqBtSEx248Cv2c6P5SQX7Dqkocxetv8JXJKyazKA586O5tV9nVKLljMQyGqw1es
W6g67MliMgeYJiZbW7a3Quob/iMweyhsiLhThkWJbdxV7VI3LEFl8z6PsvdsYu6g
HWHvonbGRobGMxVcb+YfKtMcPe33iW2dJ2IVbKKW6dZbfc4Gnw10CM4V+mFOkyA1
jmuEKXwnE54rsgd1af7Jew==
`protect END_PROTECTED
