`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J12tPgL7DDK1TLnM50u0ZFrZa+0yZp0XL5oFan30j9Rwxnb7Zf1DTRjCX4Ge0NDw
Aa27fu/KXrmFTtX/D50f0mEpr9rNtPIohsmGZh9wnzGUvgifGBD2tBcuA7Qzf+y1
1rMPlNfGs6EeTXroUbo/Yml+J6QZzpBavKB265KZB4lqGQ2wApWXPKr0VhrjMYF2
eIwvO4Z38bkUgERaepsWjrWO52tHjSuDMF5VVD+OwA58FspKto7PG+0RFt6AIBOv
aePvkmxeKvDT9XSmxLc6IijrRYzpx+Zqpj4FmoYBLXWGV8RsF7+sGIVrGmPuYsOf
QZnVCWVV4iWGKOC3HS5+0Grt6A3KFs5fNkXySWZgVJdxUCIPwJ+WgCbCKiTBLwt7
RHRjmprNr2fS9Avmt0LofsrVbDaMZyy4/4k2RNZp31jADpolhlV9OFiieCQKwOBW
ISU9s3oUK8Im1XNt1isXAnJsc8fmucR278Cc+FcodXMQ9r1FgINllpMlb7SgebPu
zsUd5hZ8wAnt5PaEAQ6iEDjjLmNVXr4DHk9kwU1Yi4CenhBVlBb3Cf3g2m8RAhzc
vBMBTPspijUsf9bvQPdi8qf9K+5nnCfDqWMwmwLZ1o7p/tWFu22AcB+yWUpEGbX0
xJBLY/v+0pg1oBXNl1thWfQs6zw+xNoufg/WKw0zw4GBz7lo5KbYey20I5xCCGl8
cRUbVHbIRUpvY0y8mVQxy+8fjvBZ+wTh2Dpu/1JPoX9Vi/bpA6SfGloMQTyNeuTD
Fes0fxDa6ZWX426JRdBJ5oZNMruB2EgzzhAA7NqD/l8C14oYXHzCfxs/s57t4eIe
V3x8XRQQwRTI3M52GBqo0RaOBbx8GdComZnPIQmMPIT4St4GIOhtSQk6XOlCxKrH
UegbFs8jtAdfcaZLHco59hQ7yTqI84Rlisj3+X+3WnB406+C24RWIIYJQdR0+9Vt
oCvWeLtrPxpVIKn4T42z7iCnGQ1MRGtsjwzsOjYUBJwVyIHba6LAmwxUoUZ0gXUd
Hhe1Dw2cgIOhOyarTALmGSP71mE766+cDYM9NXWX27AwbjOhiW9BlbI3aEk+YG9x
0yv6PK9eXFSrgWPvKAxU03+4lBUPvmkgVUw+AxO1icFUHUShLaCVbYZqW0w8d1+S
Xpbu8p5qZhmf1g1JRQRNt/J3yMTwn2af8+xQyytmN0N9w064pcHXAdQXZZPu1hCk
NNYIc1/fY+9YycKIw09JD3hTJvD5rQRbPd+E0SPpHJpL/x6V+NZsAilIjbdH5Rjs
0gSajR0NBdJHMvptYuNQrR5K5fc+zUcsRlEcPoFzYmi4v/9Xt3ExzY/6JzE/jv2D
j995B4iq/XoImaeseChBteyKeJ1t19lhhYrcbQ7mHIG2n460wRjHVI1Qrlxl2uDB
7ZoQAUfqQrXwZNiq0GWT3RLSRYnmIZSLQtAm2sY+UruUK/UBj5VhL+pNh24exBvm
Wv3MQeeKp5kt02wKikw3bE8mLVH73JgRPxguKyemAEZauuon5Q+JELncpTpPyIW7
Je3ketf0NU/xyqhHpVo4UwmdU2Cu/Juq/zTnsyCqnQRWfJR24siNK4nHCu3MYa6Q
7t7dzaMQunWzWwOq0wv25LZL3J5UN9HHTfO7wivcgJm4fqp3IcBQvTK6Ac5scAo/
clXuRAvSYorpmG3ckVF9zsVPlvxtaZ9H3P3vV32RHhvL3v/Si2ug27rdLNCLcLph
sJIa7N2U3qiVZwkwKX3VqP5P5plbKi+AOlpyz9XPjuwR+Pc2XvXBFClh0bSohOhc
dnsnT65IUC0dg3oc4rpIVda0acCq+jJsbCJEa1MDrY3pljDVINwckipLx8ZMp1/4
Yi3zfgn0eqk2FRTpVVCtAYF9XlpoQuC4dACgneeist8TZ9X03k0xhrYdzKSDDZnQ
Bh1SL21729KkAh+uDCIdBArUwHs/eetrc4S70AzpzPmJEusGZJUEAO8XYYbtiud0
GElzK5oc0letDfMMznyN0CXpuU5UUN6jFFybmXC7cTCxWwNs7f44RDqqo8E2PJxp
ltJ1lbWAx2ckXXNE2U3sokfmhzJJhxHuyeJrrv0aEYZ9Po4WoBaksxgcxYqRbHlZ
2P6BH0pF2oli1kEwjl2fOm+3J2JcGcNFBoMF9Ue34t1/CXz1TTnalj9ChP7TObWw
`protect END_PROTECTED
