`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hyi4C0TJkcmXd4A9aEI2b+/ktMhOAf5PlzEv/A0XsPls/VDUiDGXOXS+dubcWL8+
n5mguM94fS5+XJiCqwT3RfRetRsaYNhIxc7cg3WwoGpMWM512cR7bI4YHGzWMInO
TygH76AzRWQHrOpLO8Fn5KABvLDrcKFE4+SSRkrTMYdeYGX5Y/LBd8XuMOE/1tBR
PkggsJwUyFjG7FK5+2hTN0sW6dugaIUwALhiZw7i1XIRxfdGRc+2//05jjTIYaI7
XIVqhcRIJaV2eMT6S/bksF8pzOeUDpF5C8amgPduR+4VxcBi8PiocvcX3i+97Fnm
6aykbT8raUXzGPNsxQnvC5EZDYsLHSc/iYBIfpd9woX/VWDkMB4mq2acq1qpmy+T
ridFaUMAw1rP29d5wZY0WiiwfxVQ7lHYSU0aiMrrN3NW3dQx8+RK2YINyT2OH0q2
CqRV+ny1A3YR8r+T57MNpYWZ/5SIDVe0uKuhe2wri7SAG1i6YHgB7mZ7IAgp/+Z+
`protect END_PROTECTED
