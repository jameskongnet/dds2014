`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O7aagjgYeE75hR5K5yZKYZBE12L5MGl3kMoB7BwOTzdhMXhwa0t/ctnMSRT7gEzr
puKoXM+zfR7tVvC/vaNcSsdTenl0sFPD6ZWqDrSqiiveikL3WzuKx7kK9WDpLWXm
J6zx8zUjTxfaheIUr8P4+AAU+j4Xt+ddwXdAbjcZn5PrBQWCvfPLbpfqymZJkCnC
YHH4Ph4DQYG2C1IE6ATqYUEYeq786Y1rkfLPPQf1gKZ4DaBsm0n80RmMfZvucZXc
L6cFFnz2h7YUO35TgZzVP7JToijWyHvUhZQg5e+trXvZU0flDSG0l2Fv3wwNzwLz
nkl2QqmTS7WVZfcMllpV2pRuL7Oe77fUZ4zq6ge48Cui4psZl5RYdkPx7mWKjw3H
jwKrEj7/vF1Ja168/SUY/K9+cuYo2OHU4Bv/NvtsLhnEnmO4omk0fihHTwaDhDpB
FOmGXkNn0R86QZYc6YHZbBWm6iLCg6eJ+yO8R2od+yEBK+Dgg9VHpyx7UXctYiEZ
QcEXoDjuhWiOav9s2R6GC/9QEdocCu/paBymDCo5JMX4b3Vv7Rx62mFY+x4nBQJz
zHoEq81SFFeSBw9UP0oVM4otnOqfYDRMu6ZKWJm0G0fdah9SIYMbsmtV1pFu1oEd
zuKzf6KnVlVMR1LIqfUex+YN+gajON4UaI1yO2w0xwE+WFZUwUSvcDcw/kFihGkK
qwFNG2FzaQWIAOe4h6ZlimopbOIC0lJH0obiwla8dMNFgRMGZyoipST3HRfW2HVT
FAOJI+BaMnUuB3gCc81KcXxyp6BbSLQ59tA8ZjDzyTqoCLK4sukd+QGPW71ZzfwQ
IDX2/Cn09rtxVcIJmxiJfCRvJKZh0lO2hu7k4xWGUfJ9Cq+IrKBbAIrd17vjfLrN
as3sgPb2pdev/tWSn5guwU8BkNPoXv7jUiAQ4kYeQUiAIVphKMRIeP//zs63kPCo
SzaSGL0blGKhR9ULzFX2OsOQyALqSAZMfpaO/NzTnGfZ9OHs4erYxaYLjwEz4Fwh
JI3DzX+Li0eIg5STswC+6CG/vjYetzmvW1i1P0Nj2Z9jNacBv+BZY//D36bmcwOj
/WX4OwbRGe5G1BLTzkjAjP8mazGK0tpuguZDC+r3PysKKviZttreageqqrmrEPYW
r4UarRxc9gWWUMFgqu45M+er7tUy/AjZCifH9kHu+TeA2zHiSca8QFLA/v7tyjRr
o7i2xkahPXi1twwtpBWyrBAWgNIUe6Zw4jlQJ6MCRax/Rk8pgKUqMdzulXANl8qX
MsDhNWpPIOPw6ctd6ElfdCZ4NAYNHa0dEZxI+BPZwZwcuJ4HfU3e5gIjn/oSd3qN
a5ACFJ7i9yzFLmnAhRskmne3aYk31pHZvJSmLVaVL0q0x8xdBcjFoXIdNlh1SylE
rHTxL685BlSVpK1MK1z2iSVpt8Ybi0lMwI2eq9pYHMfzZctU/m06qbZ22wlsWcMC
eDApUxOFLCrp4UKXCcUmr2dmNc9T0qMKTB3qklKMeCL9sqJtUW80DH71+VNGys4C
RXiVNIq6NlPOcXNzP9TiRROtZvvbUaPkIEcbfFj4Abw1gFjL5ErQ0KSRV70Yhgo7
e+4q2kof+LZ1SnlFvZ42vde07PkEGPmpAlIWmBqOiSG4u19A35NZBXgWNqaxIVO5
z3JxAo7S2Bj5koYIkGYwlGBkr3wwHk3mrje06oWc5sxNNXA65jF8KhrIoe1TaGLg
+SrKiuJtl30x4ewNrUrtye3LPOvhskPixHr9CrKp8lGmPwQuPd+C5lcWJIX2zrpQ
3w1iadqQ67DfKEp+shWT/8EGp5wU0468hafcPXd0c6gGVgV3IYcOF4SIZGeTLYzU
PgvYeHZw3ZAEJYB2qx5XoEwDGFZva7hXzth9AmY2u8GTL7Vw7mOxbCzMC3oyRKVP
/UcJIK+J9VueFyDnpHEee+uRYbNburd2Dec5gUYoghVmgEn58EmzfnGGAZOuYxZ0
qzDNRMd+hWJue29EWodtRe2PYfbw2KumED40Y3K2NPsRHsJNQ5jYQe28a6uEUshi
KFWuKUDHs3JSUKCtyjlVlsXlidxf81Bu76pBA6Z2uluUJc3wP5G44af4Mz8bkKjf
gy0PROFQ3YdsdYR92qlVpn4DpzfuRr7uolMieXefQtr2Xm1ElHsgrN+ffVxHFoWo
R0+dZrxzkjoxpGtgZBYwgplBSVIwaN/enzGvCxGQ4Re8nPqWEXuCfDl0BCpd8lcw
86jKq8DvPAj/5+kuiIRenNvE/B+mALbJ+Dwqm++JgieTrCozIZRF2N3zPiFNRCRr
+ApWS3GbxCGTnIhsS/XEIWL0oQfvHhaac+0528ISdrfbRJnApMjnVjJ10HutB1/h
O79UL7XwQi/4zl0tLLDBSNCZAfKHJ1u2M+AxJYeFamgztuY4zH7Ph3FZ/WXBXPzU
9FsxKeSM/sXpdQ4669HgMOM9RlRgCxaDQ5sPE4qnRQhC1P+tnmyS3eb4we45cC3I
mXNEWjb+yRELBO+wnSXH+91qA9x8w4g1PuXAfUluqMuFfuDfRuXXi67WeBfCJCOj
/2TrjuYQiBEl3HnH1xkBak+6kUFpy43JUhJUPIjvRz0KLjUNk2Kgaf154FKguj//
d7ve5Oos9lhiZ7/WX0A+czYJ/7RrasfWw31+MZhXQOvmGuh95EmiIUi24ta1TQy0
qqHXZuyvXvDE3MP9UwsdFE0b69GvQnSyczLfcPLy2SbwpXN8wjoC3CFA67l+Ffpt
b2Jbc53CAHZ4TVdVJzy9dcBH4e1LnrWwG9DGqNlB3pHB4QRuQDLfteZfg4t6mkqd
a8PXZSLWvrRdjRtf07tvBzX9V3GIOYpOY/+S6ThvnQvpHZmP1BYOc8qif79dGqPa
Qd5fm/pJslc59DWSr25u/thXBMmlc/4fz7Y9UsGpVJ+m6CRuHOktALGy0mcVVrbj
tl/CynATfRpmsj44PMTRATA3cSrHBrPg/Vh+Qu0ZMWAO59qa4/XE55HCpVEP8c+t
uzCLNF9qNkVstgicZOqRuGHCx+AFh4/WRqIdMPi1qvUjL0ZAPwziAW1U1scMHd44
QGN6MiJVKE05IRPkYgeOvKxoQ385247/eZY4hDi/viMT9j21wpa/3E09/f/cbR2t
agyZ9AnnXnwQOA/cWXpjQ7uiILhpEpiZcjmX4XQGcfrnNO0BbWCA7Rg75LTFzSLX
hPD1Jd4k+U4qVOVrbeetOfm7gm5rIfBRMV3asxlgQCnrtY/O6Y4qOAiMX8qbNgMr
SxZAktkbG7lTuHpkMcrcTLr3n7pLHsOnjUTAPazuEArOeTevbpd5UYAt8bJ5CJ7w
0chGKUOfMQC2kjQL4IWxZOGdwGKX7cyEQRKEY9SOEBDT5Ygtfl3UWLY72iLeTsIK
Ln1q6vV0sRNYpcMRb8Xso2r7ESLBLLF0t4xd6/WcHu4iuo1CyjSASfKodaK6rsq2
6wVXFStMtDDO/Eh4yKpDJTTZsuGJIHnjKZyX/ajO2xpblZK8x5txMoSxlMcsmXHE
b6CO9siPjvC4NLtHhMdpgLTIDn4w3tFij820gVVlg3LdSeAVsLxQkxB6599yrH5Z
lX3uVhFbvXS0kmVQc6nLO67YylYqubHSdZdofsN+ThbmblH9+Z0MdZEVdLuCMRDh
2zv2V4ObqR65BdUH00fTcFUd6uEMH4ZqGsTi4P2A+hZzDjtfirQ7XYZiSE+AWxUI
ZBCnK8l7tcp4WWor80mb/XPNvAYFQ8sIfynqiKoz1/WyXxud51C9jbkUwlJmLZAr
eRGutyxXbzZqjLYdkNdYV4M+3sN+pP2LIrt9QwVCAXtX+IbQTQx5Y0pg6Z+7GM4q
9FKXF89vXjKbZX2csTWMj7xpBd3Od1ghB5cNC3Sxq81sr8stTtfE1R6vbMISXxOP
qk69V9phouViqFlurzct8Tuo0VW5Ut5Sn/yNalIFuZ+rKIXy8Zkm/HAc/3LEOrLf
c9dIBl7UF571JPHTXD4YnY43c0eeJVIzA2JmYh3dZ9jG1jeI/ySDBglvqQe7Jp3m
CfkZ+0pQAANNtWCXDVjauvfgNcyQA20mIi38XdvSm6rZ08PTd4/0EGKu187lx4JO
KuhEkOuZ4kDFgwG/sZ4PjBxJHu9tgod+qQaBvfeyvyLNI6mcaz+/UJ18USQ+DzQy
E7dp/mYx23r/sDZOCNVfqhPZCaROFTHHtxiGyA1autD6K5q4Em2ZhHYzXSjieDHL
MZuisaiQ9GhQ9MQsO7t7kYGpcK9QWYKW+oZu47b2NAtmO050uOwefWab8m1KTp9D
yKYDxUEi0nT//1hgsBj2vCXejspPVU42JKkgcRC75ni1d5T6H9dG3mPenFPCRP0r
mCzw8LTyZKwR51QrGmYd4uM833vxiZuCRGcsnfnpTyLL7uRbto4XUkgoudeuyeRa
VaKQDtgo1j7NAezKtQSmqj5VkKKEuQkWgQ+sWTDW0Z96TLQG6lWiyNq3U6u5a1H3
E9zWrcCC6RmFTFoOFeuxIN7nFzhi89T9xHm5QVeioLAPDhashkKOMGZ13kMoj+kG
tIyfd+MQl1cSRI0vRkZJdCNdfuL+VrB6Qa/xlICKWL0dMzMzVhuiDyx2uvs8iSvv
`protect END_PROTECTED
