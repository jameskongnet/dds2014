`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A3JOPLwUtW5im8SfMECkReqhN0ZjTbRcot9Q46+d32ywdbv71wDP1BotFxDf24h7
2x/mGzWXkI28v91DdMJG5nTbHcefgAxiGSm6IJpYQlsHEZVbPEvIF0jjresATeHN
vDPdJ/9kT+2RDV8UhuxdjB3rsBZXVQcSwBkq6cOaMtLv1cJMCX6Oa4AIKW9VOCZl
Q/I/pegPQE8Gqd/fDqVHNGX49ptyLawuDZRpyCb3ySJAoGqusc5tfzQwgBynjm7q
6dzNnMSsDxwSVyvx5fe1JagvkFi069fjeiPDEITB5E7bp0JdZ2/l3Bxf5UFwOx+f
PAAMcqXKOdAZe7DyvQ1pnMUhipJRCSP6fgwZPeCff9paRHaTaV9OAxinn0wIKj2H
FF8OR8HSfuWelPluIOUxNb2fxQ9H/mMbZkDcolpkawKFZ4yMp0yVIW+/TVu04mSq
h1iBfeDQYwjw8p1UYt0IBPH42AANXfnpsjfSLFf9aMg3sd3amYe9Vv0uLZrX2YxN
o8H3NjMvZ+Q8XxbBXnRfA5RWVeRu+jLIfl+fZTtLw2VGc8E21PPNweIxjIFrwhLu
OQziFqfAOizKxheu9zeIkA7ifTsyzpP4ip0Icu5T2JPfqpcaXa5FbwqZrIgNqg4y
eou4PdnH2TkQhX2aRkzV3hqEFTfDsi4IFuhb5c/vayw1ekuehhEvc5c0VwegGZvF
fMUFKS58NJiPzPSmY/9eXHRTCDsvGK23ngHrQ+9KMJlmJjizwvDRBuMxn/HJOTgF
PS12jvbaLEhuBYZqipr86ffhBsoxOqNAcc2IfyeO4tsRvJutfQaSQxoBaZORBK4I
/JkhfE2cX9CFClgLBKrDFc5kFN04tzeCuE1ZPkJweAVR5M9Qu+guoi/x8061sie8
VNIlmX3o00NOQKdh4O5ew3fTui35TelzSbgpInWvSXDXSV2zv9uSH+kCxomnYAW4
w1/y7CMuu/9lC3R4mss6lz2CkfFXS6tXe5uF99PZlQCWKMzyAebVUWFCTcZa2O8G
ikd5zgtiUESRd3z8ME02uTnqTFeGEjXrFjy1TKFf+p5DhDuvUS4scD9skCreUfgI
vBXTBe2aezjnl3QEz+B7FZbW7XIDoq42bmkP5AFtEU/jkiKXxLtyyiqNfSPXISXF
ySbTKMEm3pGp0ptbFWow3weiyRgMddS/1Ht5UdHfZ/kfnejzFz8EHckl6nCi9i9n
kfBbDmjXnAIEWy/+L7NLUYkPIrbkKa/K+QRi2zK2gHyhdVUAaJf17FGJjiilVB2S
phhPmZE82+GSrnfdGoSwQEL63NhYd6pz0tS72XPUkiFAEXfsO2+t13ilgxy1OiFo
Bak2tBHRCUdSCT18BCdn9CK5KYU9ErsAJgBo7YIAxHZcV4EwqHbNA/0PhqrAt1VY
WHuNs8PxDkmshEyXPdGa2EJcZYvCcXSIuEV9Zf0mbaYXUGTg+IiVNumRaxKHObit
rNA+42BQvY527uWmYtOwmp6AJ4IyGtyNnne597JaCwdskblRoKjXiv3NjQQFk99f
tttJVdTCCRfRTGi63Ns8AnblF91ZzsBbowGorcBfGbe80MOXgu1tCKEIZeUqAzZs
bWaKMY01+CjYr0WkR489HMGGL9UaRDqs2c/UXl78PgPDJmvvCnaYAYV6wI/lUUO9
AZsWf/CRwcr1qTuNDqzjhxwgXgPfjwQju7J+81mkzdFUaHxe1WdABuZZ8miuB+du
v+TAunI6IXflxoNYf0k0IG3imZmtPsB0/tbmFDcGOCx3H/K3fr7EB0xZZClaT+at
58ESLNeUxYRsQn8VykrVrac0fm8/+TgiGVQusr5+/tMbpr7aUHDgMmDwfwLSEc4O
OYAhJues/AZJbLSglI9lCYFfHjFOL1bdJEZk8eixCQab5Zd5suxW4GYXV6PuTfCn
Cgd7rOGH2lswsbaqIYdPdq5AmAghX66za+ouDP1Ikld058XSyRA98Btcz3xE0Qdm
PRhnta9rOLCi73er4M3nLPOy5nMdW/542QFoKr4q+p+p3kXmttUvFBUkLNOBd//R
xwtG4L6WkZk9QcdpQBM7alYt5htPBMdPb5mt2y6dIW5LiV9Ix8Zu1PeS2doEsn1f
aGR1Zi8+wGRdcqUV1ipN+4rMTjxqSZjlRpsl8bmrSz6tadGVtCP/leFxQ7KDTrdv
ZnPUcsuBCmzAjaq8hgjmkUmiGIPbS4thhl4cav8EYys+FB+XXL/YH22wjgQLJjRF
t5VI5MDml5ryMZGizly0VZGgzPB5IYWu5FNezPDgwiwaOGUYzcgHaC+7akus03Ag
n1BtmNu3xOAZ0DtRJUGzC5ydQQ0GuQivr1D18b6Qkupi0kaWyYsbH+neb/XhmTc4
/WZQCNvdBCC+VDdIlbXcXVwpWF2WJA6QioRJxvdG2Kpxf3dE5LtNuZQ7rCOxIJDK
M5c2eaQKkZMeN9+iLl9UhvObpRSrRhrno+S6OdeDUnRlMMkzlMOIt9tZdkenOj2p
n9t9xWHsd3Ug+weC/B33UyYkduYEsB98uvtXDN6WqLd08bp3EluG7GfK8bpUVv2H
cCKJnMj0wA45NutAPzScQrGxWJ91ie2rPXyv11XlOkQajeyC36t42YKQwTPZN+7L
J2kVYbzHXCNayw5cFTP6TPmZq9Od6tPOZFJk20EZ4h6xUi21w57uEvZeQ4mbxqbP
Qc83d3A2YgASVQo8kXGVzbWbqSxUor3qDEVtoOLBRdSuo0GJ6Oss310PqyZx9zXF
XFC+f3e+NLPZ8e5SVpQ99R+URsTr9wy+VrS/Q5vWI/3uG+QQ4Cwz9XIx/1nTPswp
fVuie0NynfypvLyFG7DPQpLZpHnveEdhuENSlQxDbA72iS418Cu9FhV8f4d4IW/4
MJyUxO6sZfZe8lRCvgTeWzXPEj74Zy+EeYuwF0CoJepAc5hayXHI+YnUiKsBBMIH
sYuXdeQ5fLn6IWwz7qPbMd1nGIHTsMnJ+MsneoxW6drW5RKgkwGaI12IEXBcA6xs
1Rja5xl+zWb9lpd7By+PODYF/x3/duadHVhsx9VBVj9bVnBNA3DUA5tCnaNBJw17
Fcy1pytCSMdvV7hi1xav5C/XxUdZMBPRrBb/Hw6hHlXso9MYgAYEdy8jQ9dBLbGP
TO5NPyPGB76UBtMlmiqGpzAjFo0BIxiy13OQ+JZE1RwSAFucwfqSShxBNh3aXr/x
nth1hk+dNPnKupID/CWVFFXapMLgGm0oeOn6KcuqYJ/ysxuugce6Mc5BQ43boN5R
BR+cE/kY3hC9Dc71puAq6qNHZXz88KGkQevR4Uu54O7LCPZF3USMgzuan5GytjCq
Qw4/TodrfiEQOJRtf05fwqMLOHw6yOCq/JjH5P/8n3f15nyM8jNUL9v/el7oH7KS
Pd2z1d0p1fFTgvq4Rbe4TWaWrUXyXzmiAUVxZy8y38/0FwKTxEKW3/Cvg396SO49
O+WeuiURJuXWWCQOhPTDaR1lLqtCcYgJysdFjW+Kduh1GSj0KsRYd3m2uzAyI+z9
h6lBygjli/5VfYYxOSRSSdT+l5VNc54vC74ILuZcmEm4PHyuXBlUocjh9WjzZRgR
boBnBZvgEkgkq4MlQhFbHNWLKD5mutIxkLHxtc9i100ZjXOs6vE5fzEFFmwjnpg2
3hFjgjgCsV/mqaOp4Jq3XpoZo40ou5DG3mPU/5OpitrkEMJNecqt9MEJPPnd5Tac
WkGPvO3fN6N3hdm4s/SNhQ9YLRlHf/raBbAW+p2UCwLLHyFfClddHnPUrT0i7KGk
w0neMLVi2XqY+ifOAY7Rv4L9NSzXb2oH2aVu/X+y1UMXBhNw8+usoyjG24j+WyXZ
Qt1Dxzt08/Ph33iMA395FeKXlxpURmLewQ1STeGSVE30mLeXhiIhx3bK51QZllJZ
Iv3Xc+dQqaUABD4L2zcD2EHCvbgJrR/EAHH6RC4CxA5sRAKh3zcC3K3wQvrjLgzq
uCJYsQWsfw6A2Lkq9V6bNi+neHhA3yJM0V7YvDMvbKmgQaCpWFZyDYC4Qd7kqmED
ZXgUbFZ+Qo8bZWvgAQuJFrw+ZGj49Z9ETGUSR5aGdAYyfh5fDmNUV2Y/3XQuOsUH
6fN3QpqZEkOo2do9Qrc8qXdqjSk+OpS27EVsjA92rhGsPQuA4sSlXjh1jQYRE9Ve
61bqevGnuunDKC/Ga/o6k3dA9mphVlNgsw/LjIRzyPrJ1Kp+erEF7h6x+0omJwux
azWXLoBcnSXX6rGieeVi+P2dcb/vfklj+JJRltx57fNsb+ftEhXpTTJ5h6d4f9/l
hSdZVGcGDnKe6mAoz5/50OiMB9bD5CoOmzmrm91E864bCZFDk0UGUswF+/EV/uLd
nrK9EsC9UNJOM5X71KeBxomEyMk57R5KVyUhKVaPNKS+Pq0LW+GZKrmVf8ZmlELr
h2pBX1S2+wL3LKmqgBQ1//5EnCS7G5XBNgp6gF1BdXizQODBAdzTljzNqxOrJhar
lfBFNzuFCBaal+1ewRhSkIhTSq6VnlwvgDGl4iASxSIvAZZJnJIakmGUgvAVHrzE
dmqap76hkvDnlJ1r2Yyi2A1FAv3itodWUae6OfiABoAL1eIZMY1XDQMfGhKsJgma
u1kf4xwG81bYt5z8j+4+zrmha0KdZDdhp7+cK6ZIKuTj0vut7Ml1K4OsxP9P5cCy
e/u8PDAHXUmxUniovHGWVcWpTkp2jF0ES5xkBaCk79+5wvuue59CEEtacVAMdniO
ailTHF6aLPE/tVjdk57YyLDK8jaHOFrmFtiCv8nQYzeE+gPVaClYSElEyreXWS6O
rbf7kuGJVcp0hjrGwWwObnSTN9/7xU8rG/VtXKpQWDFBW457TOtP0HbKlFQ6yq97
8DDYTbgnSJz97HwF2QmUWgcRey7qmQxczPHcFM0Z+BFzsCMEzwpes0QJyf9XCKRU
7WUhuhhVhXXy7Qo6O29Y22f1o5QTcAXH1QKnTpA0zjAWbpmvcloyU1xwOIZTe5l4
`protect END_PROTECTED
