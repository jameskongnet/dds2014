`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CVa0LdlY543zcNH5yb4l7ykcN4yJoRsmEtZ4+ZPW4SuNLGOTkpvBUzB96H3Yfq3I
VOmoPWFrw0twKbtBcmmw2XwDNpk5pM65uYkBavWRnIsmZ+FRQ2wSKw9BVt+pteRh
hQJ/GmZqlxrLIwZ77wAzWpADTcQRxlQt0DbaUSx+6BZkOaHMaw2PFqtZBTbqlria
5UuVWBZMWJ2XYw43uTF4RdeUfYDns4rUMTlVssyrGm19GLTGWMppOoDahtoaAZ+Z
awgDMluClCWAOYo2MskwYqcb7fKGfLRlISD6x7WHz7kj9V6QN6Q7uPhmgiLxvvB7
4oU1yGyVfmSnOgQW8OoQmVtuxxLFGcBRPGmXyvfm4we9AtpZ11jzwTrImDWta6ic
t89GlfHJOdKhrPJlgMAOZ0YGrEa1+ETv2FNI9AoV+gqeTjLe/VqAyugy5tmEQ09K
5glXHy2RhuGJt789ESp0Ng3uEyc52QaKgsLTq4K6PQZSJgteMqU+Dw4bx96jhvo8
fqAwEBstLcI4IGRWabtpAqkHRM7ThGNYbnnq0yC2iZ4YC9nfmDAxOg3pmzDRK5Da
fI3RbtWmtzcXFx1z2g7I6vq46oZ3xuoe2aj/j0QY+62g7es3HkxUDU714KE8+zNM
Wyeoao38Kixyp8Mwgb0m9TpsfDF5o26OyflJSPTvBWlDsAVEbPVSd9si5FEDJCIJ
XhdzhZGdyRBVQChoCbBxYFGHPJ2t7gcHqQXqAygvcxNYBzxrx5JsFr6o4lOxMyvP
mlEG8m7MmIh/1VkmKZN6K54XyffDrRPWJV4u68z1D87Xa3hLaSzEvr6z47t2Dwyp
bXblBV2uBJW3vUJXSuyWxF8bZZ3GxWMV85oX+/L5/V5G+p3gfKo2qK9o8aLTBUbM
OJxCbCgUQ1CuMEw+uA+L032aK1RpioxyodlOLZz/DZspc+WSs79Tb/j0ryLC7nU+
oOcjYqfPzCOQz+7hscv87UQvXFUFw9QJX+1IjzKXo/PoI4fUQYhNtI6jNpcifjfS
wR/drZGWcN5JJY2aqKl0nNWDSMAwe3lIS8JpiKLcioIGuI7OXEVSyZYI6BMkbivI
Y37nUOl/mcb5fFc6yIXysr/Jpa2rOtZo2c0GCHpcsAypio14wJnLFcUSlVVqak8M
dgot5617irfXEdIgnHlG/BwF0hJ/eAomFBnnhBCzseVqJxD6ZBcejbmgiykbNxZn
fCe1kLFkkiao+ZMm/KMALOS2Nr3yChamgiHxXXt47CQuO4OZrnGtZbI6NOdMGZxy
cvUazJTKO3Pv/qQbVs7IJuCkOb4ymRG15Uny1b4HylDAmbVYdP9grgLMDwLDye1a
wkSS2nZi4tdJ2reKFUlLqZzxxH7Zg5tbos350fE6SDQSPhGC3+wi+XpSuj6Ais6y
meicxcVLnetYmN/c/EvMValHBnxH6CDkEc3j/pzdZI3YhE0nVjOT+dUR5O8aGC2R
N32+ZRkGa4dVCIjQSfTtGJLaS8pQ9x44pT0e5W0cLE0m+cqziLE+8ltJIfjpGt7n
UQQvuMFS0x2bxXacD9yGPLVacbyiIrB77keh4BKVNZ+fZQer3sET8paU1vg384rK
hHhedos2vgyDE0tGD1VumQU6hbEVRJ55UPRH2H2DmfollZnP2CX+tCfawWUZhv9E
Iu9MpH+F4o/9NyHMMNNg/ZCozhEle2r9uwr3kRubmwNzl8QwtwI1rDpAqeNaJoX+
+tN3rkxbgXyInJLSjBDZFCNBcPIYfVSA13hF8JqdlmjO9QotaTo7rjDd20CbIHbE
t3aM3gISY9M4k06lUzIPyXUcfSYXu3LSA1DcBpe5yqQbAcaiV1QUvEOU4WcQoU6a
9idi3s1toMOLZBnJlmm1FyXHGkdnaG+JfORuhWGJOPejd+lm5p+FO0k9YDzWk/3z
qHXgESD4ZtKZXyoZOp35GC4ljx8vvfPfNR8aTd9HV3hY2aLpZxNV9A/a0TDsIetv
p3/AX5r3Ac30N+R4+wgkZ5wYqgi4r1dF2m0ZrMPReeQ4IT1owkhZ5EVaewUeSZht
o6zWdV15OHdiMn9Z2Z9ccfh/4GuO9ZJGmg2Mr7aPJ4asuooDn6k3msBxT3gYrhMt
Ee/RBiQoFuyBczNSw6DJ/M4+NTt2lhxorxxy+RUc91aC1gX+/Z48XiGAPgqkUeJB
uT7NxaHvFRZItmG44rTdqBbFpTCUxi5/0I3bkx9dYZr37KqiUv73j1+hzc+x7P/S
717lNGKXUSBGld4ZvCsBVY1BOP1CrZMVxzTFxnGSPyk8qwM4cM7+f8PbOuyKj725
Fvh9pAlOTjki30Vr0DDjoY4wD2H1/6yWMF2VrmFAfN2optyr0OgeO8prxmKql8f4
QDVnmgdzj99Tgv+dte3vfNHE1TKrPjQCE51ESgfp9pyiiXzqabNt/EhOM1YUqb4A
CvvPMnr0b2GOKoOxsxtgc4/D66eqIDHcRVLfnGyrWQCXYirvCMRCtH6PoIF6NWLZ
BDHHT+S1Z0MGP6QnNXi+hF+rLbndwVFNSCTTzi1tzE/dhhOkril/pbtN7jKIYf9G
56zDg7R178te5EXrD9NpLdXJrLVMcIKJ+UvCsh66Ql3waeHzprx2Uq2Ji15QkQIf
NlcpI0LwNc6eIlpiano91Ie6fQsng+Vg9YpuDJfiCUQo9UaZtbJeL6bKD+SABAbs
vE5B0Pn00t0xEQRZ0B/DaPM6IszNQyoSTuPT4izT8wRLvyt2IDgfbRnWETb6ZHn5
Vmn6Y9opoYhqmP1MYpZ8rLh0E0T+d9hIsK8NUlhfb1ewrKsDOoqmr5cQ0sNwjuhq
RFqfboqTXYA36EpkD4pSSNB7BGw188T8j1KjEEBuOsfChaaxlYRukjwVJXJBiDzw
Ay302LP0ZSsJeANJeId7j7+gehFnNhdGHGKmM8dpDYsn9tyA/dyhNHcbnJa4lkdP
dF/bpmJFe8gnVZnMmFYZjEN6mwG/6Mw2qXpa1Xq2N26Oh/830bw+kR0w8zxOpDwJ
jGFpNs8HUBRkoN1gdbYQtHU34RwSk8sxVoMrBipxJkTuYdyZ3YfYNRUKJxtjRYJh
M5uZ52xZhYCPGSY22TEa++wHslhV41ThhVJYnWfTXSSdMjNMxeORdHn+wcc4SkpY
G1mhOTjlCR2Qy0HW6SdXa+1FCAivGk2Lpdb/vyl7KVpZuU2t+MQxBScQmDaDK9AH
l5Axa+acvAvR9jnBaLIshqQfom9SsTgELdHJkkpDHaSqc2AHSuGRNLLY3H9j+2FA
t9mfqhLVnLHZQxcWY8skxdGhIsBIWNd0nZAgkbUG2TTt5m17DQf3nsm4xraoUSIh
G8Kf85GxehxwKkGrZgljsvUz32NfdvYUfCeShspFXIo0NYkKd5g0/JZT0xvaw32K
bGb57EPyteUkGA5OD0I3x87Nt8IIV29ZQeI2SFoRhG86T9RNolftN9PwHFX20Pq+
8j9q120R8xXkj/ItWMNy2Cd2KZJcJxwqIcJd/gUz6tNFD21vNWHlRL1C/bX7OFdr
56CxFfAnxp/ae9GkmK8Z7+h/BC2t6fwpMdmZHZCNwOho5t8t7weKTHhO1Iu7ZXnQ
lh0zaUxHURdoFLchJVfVYe/sCmp3QOMAVvH2Tx6VgUO19+kosRgp31mU1UU6EiWD
E6h0ucG2cSNkQhI0xv3egF1CDBxIPFTQr3Sa0dM0LIJ/cV6dxAoNqV5OT8qicS7l
Ms/dQMpVPDDumekWTgEcWdpGcFdYZp4oT8X3eUiwI+SRuR2qi0SVlq4YU44osfiO
LoVZYg7/93++KC9Q+d79M8E56789bRe5gs+RtK3csNl1MChn8yL5MaRX7F77wd0A
wdBRKWoD/c5LdTd8ab+8dQKa2s2z+R6MW05fE2FRdLE0QlluIuR/QrhZFpj6b6Mx
VQmK03rz+dmlRTG44dnnbeTEsa45TbuBBEurY/0477/7/GtZJViCPdA8G5VDIlD0
U9TyVfdeahftwP/qyzV8TiRgJbQWqKJQat8ywPMvTLEAXVtFCOMDT6oRSzgF3VsK
0nSAbI81Ro/dv2iC1V/evrRcHgCZXmtty5NPVG8VbpF3IEUb7BMTw+H+yafo/Kqs
F5b/juwPrvvK9KiDkNLgN/opQVoRabHt4aIgkOtgHU8h2c5TAkwulR8obitMhkX4
DHeUC+vgmU+F9HvYH/bNz0NCQXM9zXq6+b6r7aF2pkKfq+aadmgG+SOJs9nf/BRf
ApUcupe/tXV8/7kAno4erI2jO+PgQSkxgP+yHdv/ujf8/o+zjdI4Edpj3aMYt2RN
R0lkK6BmcA32zsiYU3HJDfOVFJNHriPdfviuQ09OVcb5V/awMJvtX0Kz9ORULnEj
35EInTXNX/q6UCRhUVp0mZAG74UqCxCesZkfaP7Hy5wMPXen/AP9BXbYW5WF7K9i
HU5y/DwA469G1/Gj6pAT6r0bxEtfFWiu7o6LIsX9M5kfgNxiDrAt38TmMMWac29B
`protect END_PROTECTED
