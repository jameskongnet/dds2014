`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K8oOgD4cda93JastQrwCHb3NjaGhLT6LOus6g1ZCozMLpAKaiI5C66ErXbZsvtT3
Q3wrZ4BS0Sk46woOUKhrQ+7V0ZyjlZxvWqjhs6Fd84TXwPM7R/bD8FRi5ZbzkEdf
xPPt1w/kEXmuadrlj1jbmMFa3Jx27DLM7gwyEMit7a/HL5efp4ZEsYu0ZMuDJEqN
klvp04vrTzcQJ4xRSD04lJvTBUB9Qtwllz2i63j+hamE9zIXiv1j7T/+1CnMcYib
MMVj7QVKU9Rw6D5oRlu6qy5PKr4Zeg0Ffe1RYkSrQHYk3lAuTs7nZLaQZChXMfWc
8HURFDHdHmRHhPHFMTQ9zQIFpICz8iXbeA8NeSc//8v4uI5JpIxA3OQpleI2ZHtc
sBs5sxBQ4azMzBxgYsuGV8IxiQTO5T79x/XwecmoOVyseDbs3dNWlDbnCKAiUMHs
vPbRCOk+791hOPsE7XOhL1Xeb73t9udriPcJq6aSFARg2QtJPHDw/OYQN922jRoX
`protect END_PROTECTED
