`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9L5eaQRw/zs96iKt55bnWEEpuOnPrid8LM/dmo6dQ3XEa/GmeRYM8d2Rq9VbjE2
ZnMSKFgEpAsNfU/i/RXJb5fLoKhUtzElAX0H697Ub/N9WRks+e0T1DClA9afSkgx
FOwi4zoCi6qJTCMG5lFnxA3d6thdKtEBhuZJznZTqf2UMYxdHP72rhHZKf3AElFy
roe07zvUiUyqnSbebTgqd1axXRA21u2JVslvT8MYeRsxGrdeodXJ7waAkVeBDf6V
rfptvKRwlijEUeAkClJyTKopB2843rstiIuYKnq8Nhm6u3v7Ib/TgtfLx7i6lpTG
pX8TZkZleWFGs5/VOjsItRYBjIMuhRuDRbQhHmGZ8g0pjvHN2RAM6HOamscWKRET
BBPmacGIX98fTKYGLLx6S7+8+ih3PMflneqsYBIG5NnRyfMMKdb3+AHcFKIzQMXP
+7HXPh3Me9PS4nbiwHfZU2Npj1Ofk74p0ppALbq2pBVZ3GjFRMg7jdP6UwkTQjV9
rUAiHTbLnJ6lqSvi/A4iUqKMT/4kWw9aWluBQZV7zqcLmonZR4UWBAR5iTMtJE+t
4ZVSdhgvl40pO1aXDVPn2D4IvHd1pCWtAmPklW9F3tOwDF0VRhZba8RwKPcz564Y
3G5jVPnmpLOC6MJ6Jd5icea19h/pm/U1jrAmT/3Ez+AeLoILj8ROGzepgwl2JzYt
VuqR1mb+QIsL137WeC66YMjDxsckyWbsAVwk7U7NHJu/s06kNY1fsCTm1nv3aYzW
z15dX2FXOgN60tZ66ut9JQ/toeXMv9CEMhwMwzkfH5w/nx5VeyvJQE1WDir+U3nr
ZXm5RflyE7UaVkaA4hYiTW16aFC8tOIr5Bh/eKg4cdY70/ldqFaLTnqSyxAsLcEx
Rrw25iFRSgx/BJBbrLm/lOFUNpmXabzx5+emvrs1uTbIwz0tZcch378Cyx8ypkMs
ccu7wdvnAHSyZntgPt0WMPqrN5Asa8m8jZcaNtfM//R1NaEdKq6t9TiUCNWpJTti
ZlGC2PNwcMVZzhdduE/BfiVh2WvaZiPLcr4a3Y2AIUrn+16hs2XDbZ35DnBR6MhO
ly19gMeMCXuBFwiw9EeK64uJWNkjkC8v5iuv+MNFoth4CPQx7lJ8lOsa4c8USP0F
qp6WdBU66xLH/WeQTzctWLLYdB+6a3VUtroheErppdKQwoJGXDh2IJEI4CthATEQ
R3PR9NwyEytcUh7/yUR0rbhwLoVWSXKf/fRDVmyEGEZxvQ6HhFAHGM6NQrQjLGFU
ES5ZrRssHN1TNvwo0JQVbw6B7c/lf3gUaJyHIFbQryboj/Rtw9NNfcn+xIRPF6Sb
B93wZj1cVLbsst8GoPldVLid+htyTqbWDXyjEWXwZF4iOlg4qWj8lylqvExnYew8
s7T82skoneokG2ruB/rfnrTYkMexBW1acCv6lD2+w9vWLjNh7x6C04VsOM835Evf
eBO0oXYSZLw2w/khnh5OtvY5Nmpf3fYfjC3c+20eYtC3jcJpopHUrhyDr2ftoZtu
YTH1j7Y0MFEeZPtbhdMSvpNXRb0BPfTvnp2DcmCqk701tgnqJ/IL9583bpvEWo/5
Kp8T1I7VFD/5Gd7p5erLnvkmYiPz6hoSAY8YtOogwcu76+ZIao1rFVf0FmH4Wf9A
FgO53T4MYu9rZ/JFOwvR0Um8OM4VaUui0ShoJbXzjydNYQ0w+pvSqFFZbPJNxa68
Bbnz6CbPnVW+EqshD75vUP4noGpi5NITCCXoGZMO+uVR/ACel/dO3oMPwAcC0jGP
ka2hAFL4mjCmgncOAgE2G6boABZ61lWNa+l/AEyW/OqfUvGY3Zl/96ERcT+Jujqv
QmJKbqHBmSArcGHZj+WvsW+Rfy5U8AGS9fyUxiDw7jd7RKa/ItoYEQ+ZYxtf+IBH
u9VOm/hWkXz3GygGvkuz+jTfi8gGuxhT95d6BJiTZr/Nt32QJB+MhWVHWwqGVHPp
C3eQ/l1vE9RkFhaVJXbZ1wjXoxBbLah7qcLn5q5Q0q4UEmFTvRbXZJ6+OuGOIimd
oRmtcOCyO+9fQUaFLILfbYR55IIe6gWyftXXZXd0QR2vURW/yel5G5vp+TGcLZn2
yCgs3K073Q0tFE+eKc+3mErv+5ojyd4vAJD6wAwvlDyPpkfgp3TdtbcZta/Y+9Md
HJZt97Lt0XniUIDrOWULIzS4oClIYuVpvWD54xMAtO0thy+IOzgayRerXqcBb4Hq
3xWkHlVZGjo3U5WX97eZ0CqxdBDHsEgQ5dwSbp8siq0HrqWOwbWU2Y9e8VFEq45S
VMnJnfJZskr+j5NmQtV8M1pQJkYi+DTjLpMi+VxxN+FR930DwiuIXG0XZXhChHA9
JW5PquIJsWCg09HoIZb56AEEpq0Y3g0LBgrhK7F5lNMUwDCQ5Tge37XU7YPX0jtX
3Sz9aLUgsxBMbNp+qqGa5E1JXawgnbpHs3Et0pjbCbso3BncMKofNTmMGp1954Dx
f5cGNQpqLA7GvCEy9BK0mcRHA4ZmayuBEmKnCDw/PtiEtMwpwSJq+rUtpkNmoL1z
/yix4gtxh+FIgmK5Ek+OLQ3rLmBVi82txT2Bk+zVLwvHfnfpE9HU8omq1wFWde64
8qHB0qmD7xmMmj7C5EB6OTXYvyuO9qRLx/Js8a9xMyUlBBe2cytJjbJ0HEMs8t99
K13edHO/uE9XQ7R9VyCJLU0jI0/m4W2h3ofITEvoRtctfr4K9/RIg2mk5bLUTXeb
PRcnL4GuryTL+193ZFVi3r2rBFfCL+gWIiMZjq8IBmfaXhOixScHSXLRiP6ljeth
1fbZSIzoc6Mr7jYoS2HJ0rEVrcUjLzXpNzUEMcLy8ihsM6F2RfT2eiO96jEfLKUY
r0qsgDpHpqeim9aLwbAC4BzviqWKj8VHKUjOCAQE/XqYKZL1ahNOio//Q/KUiYcm
PobDbFYmNBU6Plplj1b55mtJChdIbraA637SSh/IdPAJKsdZB6ZO3MGnmxcRYxmo
DRxxNzZFCQn6IDcu5Z8Q0ZmWpi7QH1jiDT+GWhiSM9+AFKZnDu1gbIxVgnS8PxXq
WwU+luOr1QLcagROJrBoTEoCerABBLNGsXHCSZm0lA3kJdmsU6jrKhqDNwYQubQ5
JSxSB+kGaFrvCz1hioKCn3Vp394kj6IgzDA7Grsm/Gd9e7qE+uHgqxeFqMQ4Uj7O
vuNR0ivFmBbam78gY6sDs1F0icsRY7wi3536McCbYrkaJpG7b++zXsH2CUS5o5iD
h0GUqj+DqWyp6B0ZMNmQRXZJ5o/CUivm67KpXO1OnnxELf1qgTE9UniRW4Vh3GKQ
cwWNxmxtlvzDFygY6XqMEDaVnoyyqYPFsBmrGF25gxX5nQpen82gwVdNxBNZj4ig
7c1ywg10jDWc70sFog9hvpNaQQuQWBV+GNfS8IzuoxBzFANxMlgePXNwEfhOmZzn
XAZZ8zr+Eq4m3aLDqnhEBrFhJLk6jj6iUotnnIXlwONu6naH3OKbqnfHZECPiQL8
FP6NAa3QOW941exkIC85io+bzQVQlhKQO/3lOglsnYbXguniZ7XMOb0mZwbBQSqx
qDRPhAySbyZEJfwmZpX8z7WLeOvPupPJSAyMP5x8C3NA45DpVpbmP96WVf+RcyvD
5QAzblf0tmN0FmwqYMlt1Q+cI3NRoU7O9yir6SoYIDXh+1i3qHuT6YKtZp2J59Dm
FG381Vwj3iloL7I0J/Mp42v9yNCtf4KAXpOTEzw9mwVkuadj0b4MsFkxWzRYANiC
+czStMuMv8RI0uJf/+wAUjrnj58yS4c9fbBl5lVIPJhQcnOnrFfWBO6w5xx6TYfi
9svQ862qxhyYIU8iMl7jxbIAiuIL8SbQ1Snnjr8+YR8aSgmfaMz9upTqJffJ89AX
HrbPXIaqnOOK+fH4ArrkAU4OfW59njzjLJExG3wCyrgjYq4jd+rCsRkEwu+al8OG
xJWqGHNAW2Gb3QsdUrLTMGIfecMl1U43ziqTj/g9GdGemYmQ9b4JfWDLEOx7rrcM
JkG4UHCLhxU2tDHp/BaHGoz91EeWhrpTBB55XOjL3jM4caer0eKUaOu5R5JC0Uju
wdmRfZ3pgsAryXCLoaRew6YXiss52MPEuVWbNuboKlB/TYsPKRTFo3IjetYNa5EN
I2cbI5zbHSci5thl7Uq/gzOIdK2zl0Fg3JU21k8N3hr78w+VGoGBVs2eEfvqRfsM
XOo2KfuOwtMx73qII4S0g/YNRQKOIdTh6bDRwfNnnA9XBVYo+dXVD0sGvNM+rnq+
x1goduQtx1+/ZdRTvEyU1pe0s8hoxgpeoC6mv0RcNh7Fl0Zb77GQtPkM748SFk9y
ABM3C+Lp+/eW5BImS8oXocSKDOHNoxNI3xk8E5Scf5uCHApzxDM/UqLDR4tI6Tkn
CF+5YhsxhdXj12VAMJ9FwE5EXQwNyzADvXwHgnLGtn5cnUtO8gj918Bg+KudFXS1
VVuGe1VOmpG3EODlX3wm4pVE5MSlug0bfPLrMVKBeKvId12sfSECoiNPLGd24ZGr
UXX4bzX3NZOxenPPxHS1N4VVSVYkQqc4xkq6IuIIvI0K0AeT9qnYP8KcUrTJqfaY
wmpZg3aYoiM78nXLU3d4EuPgH/Nd9REDYtGVKQTfkY+1uurA3eaDxBECYmrvYceX
V+Y9ZMw4LX0qiVBkUE5O9sN8g6atxq8WCOq7hBxeYrCYkzu6mxVI+dTScYpL1Q83
4SuGseNG/5vpHZgTegjCb31TT4/ygtvea8atc9JFh8E0mZ3eIiy66MKoVjp551o7
1sKxO9NqhvpadSS8a617VsqFQFUzo5muExa6PGQS36exmI0OqzZrJkn4RK4A6qIs
kx0Y0bkNJgQZ1E3A0JgBjeAzm95J+mPHcaVovJQtmtDXIM/kLD66T3relJ1/K94f
PdjyzIb6XvZVKIVT/lndIa5IycptC/6h2uL9Pmk5PhY21dKGKngUqo2W1qrdfr9a
O/KO6F8vYBOD9jPJ+9fzz4/gfgPhxAPdAr6hq4ok6ypH5e3MEfs0pm1ymBTxpfY+
sO5EIU7d0EfV+J4GSr0CoMgrQDBPGE6S/xybGfUl2kf4Tf6rEA1ymGEOjul02cfc
MHu6+O6HUdyjQIRGu15EQervH+4i6C2BD0F+S+t+5kAkCE+rRgRzm6eGoQ4iPqkA
pqKjpNu3mkiRwzoStAP2eKht+7GegHAccwEWidcDbblaLV+ZjOwDN4FvR0PW3NkO
c7oR0KznzNMIEZqrZI62v77IesYmk/DA39abZ6IzY2klwZWlq1VDikKIaHt27DdK
TCReLkosCRHDVlAc0RmvNujQlT7VqPCFPs6Z4Ln+EXeAtt2BdxdKwRAUbMCnJsme
3byqK0PnahsEYGKjl+3/RpHrkdNSlH1UFpTzduyWjkmeMzqtcuejPc1im0PkedYB
wQ5AWvylYnq+szyAasvWkj4Ax45v2cPZiuHRspJCOFCwvvYTgxPfN6MDpoIW9BiC
HZpB9fgeDmL3Z5N6TjtYS/oaaztn1SHwH+/WBxguam5iCvk/8QS99OFf98p90Nq0
h8yL60YyW/G4jq3Ayx7QRZIn9/5189gQQNHJ9x3ERZ6+QRuCe3dhg82mLpHee5n5
UemsybmL4KHIht96qjbqunqP6gb5omyKRk5d+ouarBkf8KGE3YjwIxytTE3Q9ceT
S2oIcGVUWmZZXn6CI7m69af/zEk/ULzWlrQLgw6CcS3YkhCMR07jrMqBb9zkfoyK
R2D1gHfJCT2qczI6nBvZJMe363vQ4vzR4UKUo+r3B9sbHxf57ggNewxO1ksfX4Qy
XsLmIAX0WsYfIMyZWte2WBY4oxFi2/M/hCLOlBTlXDooL/vmT9SFoxJigv/Z0NeX
Tborxt/fMiVCpoSMAiKD9WZFN4RmQ6pahvdX1WJw95Zcd4my0Eyopi2/2fE3ONgQ
W9er+8VveTzaCxh9ovLE7EJVIXTuVvFXX3exs9NUsHWZwEIrrhHw6MvsOGynGso6
MFmToJXLMozsDrARmUZD69zF2kGv896LZx2pqkqk7F4zY8fktNqgsWG42aJRnfTB
Y1Ve4j9wvb1+5OqRs+YUt7udwCGdjFadN4764wycFR2jkF/YYPnL/ojLxE/Q7WIQ
ViaDzBe2GzS3n4R5Zy1/+D4vDuAa8TWwzfWmZNYs0zJJOBPp0koDM/uJs/WaatpT
Jc6pEpY5ii0f8AV5DNFLEzHnvNPdu6Mg/JRIKWyNuP2SYJBK49p1ieEVAyKl9kNC
Ke3uR8MHimzyRBKbus60yUbDZFVzQT72QovXrgMiU1te8jZPnrMDUrGOqokyOYvU
VqtvPqWbCWSUObKWOLl+p0RFTLKNcxCvAMwUXSrehce9ugQRwjg3nelPHf8V5FgX
eOcH6sJ8pJGxzCIviuF4ZTiPHqxYzKGO6XjUqjKuzgnFHe21a1ataIfcX1/MlL6i
Wx7ZTaixS9j0Ona9pR5P47cipnD9kfl5inS71AU8rMn3PfLK4Vo13HYJrjXlCUcv
06lEsesRLOqZ+wrI83XFZ094G9Axmhk5rkfUPCap4jra530TP/MNSyQTc/4iLDJa
2Ba0fOiECkgbYYwUggGmVBUB/ynezpcXk+K1IrFWSsoyWNmdr1YBDFQFHYC01b+f
ZHrn7/4meNy8jL0ufbP7fBy5KgzrEEXDiHCFEZEmPcZy7BpUWadlcX5AjDk6WJaS
yqkjmBJmo1X8hAh6+Efmf577J/O1ImTm+GSvojFmWMxomC+DDsLYHG1GTBhMpmz4
iEFu/xGk9MR+jmhLfDNFRkx9ltLr2pEtJlG7MMjIxttIl/dTik15TCmP4zJ+yaTo
hxQ3YNS84emvRJct1rF51AEqvhT7HPjgcR45goAsyC60ijI+N0Nar/U4QdLFMXXx
UP7HE5l4fUUiSMsT/RI4VEtGcs82EcRztWahsD9ujUlPuqLId8ge+lMZnyEJNcNJ
Sd+ZezGlPWYB93ce95NC4nyY/LKjH3gdWU4bj9l2OAuwEOv10l379bQF4ZJQ+gFu
KTonJhXvjYsVY2BsiT3IEa7bKMIKndcJeunsw1ojD24XK9w+VfBmErJM7VDxzfNU
iLzGyfS//yR5NfvOTFIAygydgcWPRFW7OEGvbCxkVg8/f4irvhxqKXSW72gLysav
ub/oFXng4OvtoCaxkUcCBpubI5yXuECqioEAfUY1Y+RIWQtWBQTdRX3og15l+NNB
bH9LED9F3X4ea2jFU/hw+Z60a6TaiJ1ckXYNL2q5Ib3LSixYIMraUiHrGbMvoJWJ
TMbObTb3ha1Awd4djqg4uZnGOtWLFqrE4bidMeAvb4k7Am/oOWFcil5GP/9lwdFo
RbmREBJNxBMfQnKKnpvrfADh+1YSwgOq+rZhc7lIOghOKD5GqUIKjlLfqeOhPhZ7
MVlTFJti6czYpvu5pBBEmuuD2XFS66qZnvHHYPqtCbuktX1sgL1Xb6l6oBk4Wuxo
kaPUEKSoURFe42RoMrsMxlWuYBMt0zMEN3PpIrsufiqXaipDLyr9/oGNiJlAa3W1
Nu92g2PCDTAlTfFwRi9f32o20n1jddaq0D0SCeduppK+EpI639gQkDYfqnAZDE//
ErUeNlvMXlb3dPxsBOUyIRsGKpXAehxXMpSXnLGztBrNWXV3LaCiHWHP8Wg6GJUR
5QArwGUgyv+g1ZHQjBzGqLY/LSG5oHd1NeeTpm3qg8fMzQ0j08dxsOxr+W+J78Zm
h9jzz6XQE0ksF0aGhMix9mGCDQQnIHA+uFaKhp/N2fohbrrDKCLtXN/IKngePm0m
OoH77klHpfpNMxJgTsPdsb/3e7MHY1LIfSWHs8cCoIRTTsRobCj4EDbcvqDTiBIa
RrgkQHhBfg5toGCcsZsELNRBMO4jIhg8nJsoICDmAJFHnZDS3DbX941fndK0ZtKc
HOzWG45QyM0PMQIIYu5Wt4fUVqk9PDb5/2LjA2bBSL1mTZnmgNpOx+nEa5388rtq
VlQcdaf+7SQt5AloQDlfku6vCZncTH1Q7Kdlt97CImFmmC8w3NJEHRt+y+PBLaUX
+tO5dqrvnwhTni7xQbI35UNhpTy9ZnJ1KFBa29oRsUejQVg6GsDxYfxTldcyUWGY
qz0wGWMOCDH9P4cg4uC7T9JxCLRffcp6/foeRK4QvJAC0LxYgSMJYEsMn7MYgum0
HhTkEtvZ2AbJi1tSRANkbZsqLy3jL4tcQhgQne+AkULMI31GKV5K0PUezLYWAq5M
p9kZ8ru2zct0kkOGBIhXapekv/FR/ra+BTRjSC2WaxujjSPOdvhCksLpAx3wpy9d
Bfkn1avYxCdbApObeYXhWVwWu9VHG9a8mo+bCsFEmt6hK6lb27zu/9GgTbx4V3Qu
kk4jFl7Cixt6G+6TufnIUpRV703lTzH5rzTSSgL67a8imQqlufN9o71yR+T00B4Y
njG74hiuoD9Se9aZ9CSB9dLi0yfh0Rilg5ocBqVnqG/zpZ+J6+WPRD+8jIX7jb3K
rERKNxh6HmF4SSX+O6KA4lZVGyadFSysxLyo0YkRFNeMZ2NrTWM2MIrbJFfn1X7J
Mt/j0elJluWhPMasLfEeE14ZOL2Wg2UMOO3/XWFbsbTiZIFdtfOw+3YU5aaj7n8E
jLCqGeKWrwkFhE2PqV7QCFh9h43uCGzWMhGDbPSMcK0722wrQ3OCOwaoFkbAL71g
718ihEe7h6Ub1Z5v/+KomhtrJrPQJ+fMuUpH9bFN3qNKZGZ2qJYIT8Exb5A2OjOA
c7CFjLRVmbh7YlAX+hJ7O0R/3On/ooNAyo+aZFQbeUCRwKo6LX5twS3bgTt8oEfD
BrVrx74SBX6SLb/2qRxwChxN0Z5xraXBSg6ja/3sYnUb2QA9NKt+OIU5cX/tSHTg
KNhhlUOGlzILvFme37e9yRs8/4GPuYHTPTSZlm/MezEgCkVO5C+7T2x93FJmpVcu
Dd1EtV63luuuwJgK40nc3j5QO3SgtOLX+ECRJ50YelhXzGPvXZURPIeCWCZ/ljtz
w1ln+qkGv4SH28N44EuuHRDs/63lH2QaEh+yy6FWgp9xpB061WKya96eBCV147Gw
sKlUJJkAksFq2ri5j9X0VqfSu0y2h4rOB1etX4zkD1RJfBrymQ1mKzzoXFx8LmZk
NGmlQXKpX7izNYDrExPvoj60eq0YawBEdyJZNs/SwBtVxzOKwYjE2GcKMkXibL6u
SdLWP0RkvnCfLAxKPfVmHIKMCSyx5doNiU20mb7UVIogBtERkGjcM5Kv2jwZT2qp
FcJJtWfjG25amczjhWOXl4Dk/ssw9J6cp5y9Eo6xzpzvyAdr7krUwqv8Q9appUWv
ITwABlrEcrx5YjwcS8iT3MqfS32lUihr9h2ADA4pjbpPUskzBcKyda312VF2er7b
w1aQcR8qVjhY6NmKEgAWmUm8H3mmfAQ88ET1Jq+a0weC6NAo5cUaeujQJk5XGBEW
4xD8ZiWNkjpOeND2tH+wR3Jz+7pLiiz74q/q2gzOV7/pNs+wjQ7lmOJ58Q6pfD1u
RlkzP8idHEC75jFGmwbGPQ==
`protect END_PROTECTED
