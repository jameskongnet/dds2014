`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hsvWpSb1Vde8peoC2dBp+nfykmGo2awkE2jJ7XGDQRlgYdGDK72VSVHJVrXSJzwa
RbH3Ogk92JaF1gCELHDGy7LZILFaDQ9iz1b0wZ7Z50kCpCs+2tpj7fEQU74BX0SP
P00vVGje45+j+NsPHlh7izqNLXuDRu3OtnUN9fdtJwvmLCPLr1d029GhpQTePJz3
AZyYTdr3mhH626h7mL7vM0B5HmsucbBrX+dXT2LTLvpIjTR0z1DMMz7QsLXjF2ZT
9FjO34tR1tRNERZLh4Gvc+AkVlKJOvxg9RzKArFi20x81rHtCVT/1+JVYeiOALV6
OP64RFhF/Y5alUMht9Pno9YF+gbIgqqMn6Lu7IGpEyyAzQbmy1r6YuSMsY/FBTJr
FzY1bKSmWLWgzBl6fktnr1V56Yk15euW5UUsD9mXRUtCqkOwhcgDLRQftm1ZERbw
svSAciQbnW1VoZEJP7A+DQv13XgDJvvf4n2OSYPRbhgZ9AH4DxmDOV/h4uQrhAs4
S7JKZpGCcCwBp/IZLCGo6sOts8Nr04UUVIUu0br72PD5gdE6qv9GkcuUwFCW6/3e
5JXr0kShinpSU0T6dyENBlccx4XE5qSxOJrEcSOu6LvEuNGEzOc7dkZDjhAjENWR
Hi0o0fWZoRrlcZ7Wnx8uhJh29MGstltUaQw5dAGXrSs7VQ65AfRdZAskK4JGt6Vo
3FqrDQtBSd9LcnB1lbtk0eBjHtVouJjGE+OnC2kSPrm24lJ5PzJL758de4eU3vWI
Z3LfpIwHSYaxvSoUHGnBQkZoYfByux2yA99xh6/1Drv9cAhB9fiwEZmhPIjHik/G
lN52ensbLTEC4NsCePgT0RB2a9+3P6vtUtEsDHkr74jt/zlIW2Z2RmW5NeIIvXyh
0P8Rj3hH0Ngjlgc2eWcmS/dSPdt1y4rNeCbyaoLDnRipK82bednlgAgn0tH6sriW
hMqg98AMIi2chaQkUebaoOD00JafHrTG+VWw3F4OYVU4bgt7cTg3xO1vXMVMR4eh
FR+ZFiRNn7icK/eUXKZ141VBvKGKJY8CvnTMWeZFqrGmp9CoHCH88ohpWgE9kB/J
MB0IKxEqgzfGZUx/4QQ9m52a5mZOnXuuQtueWUorabrBitvmtw2roqCdA3rDsML6
7r/ayQ0y+0lLq6dxTggjSpt5pInI0lJKH6r3xSL2SJyV3tceyol0NImXobrcqFrj
8WSeUMWK9RAtIoVfx2KIombk+040F25qXPCA/D+2iBYa3lRxyhomgvCZklpe2kih
`protect END_PROTECTED
