`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fG9qgO/bwSYXia/B+Z/eIEeit74lWY+H0eSB5RfPiVNAcbAXdGuWCcJlS4ZzG5H6
cODQyRFlpbo3Q5jTOTtrGwJIeCl/8hhp7PgSFZUM9CHkXxDJWcExHroeGHBaICkM
wy4k86M9Fn5tAJ1kySNswrkzJ/rvwtRmmlfCLdOr7VE6YFgunIP90aqwnR8CoFfe
/NIZ33i+50Sum2yDkN0fpAKLSyKAtzbKmy2OV+LZLuWXZ81EBTcFgHrTSRN/J7k/
K3rLzoxvxT9p3ruQG4cqAR10Yrjf36IyUzRpc+D/u9hEM+MKbSl9KME93Rra+ViY
B/z8SuIRQKEhjFv5oH+DqONWMo5heyB1hVwmhGgtTbHhaMVD7aUrKE+YK+wGG+o/
6sqYMtMe7tw24laUyR9ZvEPsLhskUOSpe0Hz2T25DkL9B+VElUp1VP9bYY3A7els
7/nlxj8NcUPn/YTvX2T2AmtLOas2fSaQy9xpCjuJRUvLbMveHRPLakgefu7XMnY/
NHJlAjr7kUVM9dh/QzpHdjenk55PdFXE7k+/CGHQniJe9v8pLfvt1LGALexIYaKc
gQ+ZEC42PSKwPhLlV+m2/G0CGfsRqYxq9/JGbZtbQLhJmmATWJXbz7lQCl2wxlFO
aNTc2bgKosm5iHPjiUuUst8UdBbIQ7Hpos45j4EAHYQs0iQj6QhCps4z0nD23nDJ
3UBDPGHzLYuFtkNtLZVjsuaQxkuu/xYFm2fwAimrCHcBvkKL7c4eQv0SpWwapmc2
L1WittXH4YpinFQ5QABCacRx6iQiaBGqnRAO9B/b53QwHvXPPq3Tj+/kT8Kt3Dhs
fQeQwQLVEUQEfr1C0G8q7+R6VDSJHRSge+BNDy6P5rdKOUKa6TSDgQsBhXeLEfNR
412csSJ6cAE6VEVB+SMEeC/Ld/FuZlBVLqVY1J75Mblfw8qtAZq4quryCYLzfurD
u0H4mpZqY6j48W/3A/TcVHEqWGNoCX/eu9H2EoLrq32xV2zEdcYJUVMbZFUR1a24
HzjLs0FiWlDJKTLG+dVg8angbL1wwnV1r0wcWdPrRIeR+Rw0D6NA20vXqVBVBZGw
Fu9VQav0wJjpNK4Q2s06ucgQX69NmxDx/qGaQ+//YmTos51vbk3B6ykISk5rwTcu
OCxxD7waDWGFkB+hmtkEvV+K9AAFg96+fRHjMbg7o10tA43UScHSGN6avpPy9nsA
dUIIEbtZ9J0vaqCHSy4xVHE/hF6wIr3N1yQQxQsgVDueG7lEsGiynQCclzesIPe+
8pU2nw1SrpZl2b3lgO/GrfyBFH8yo9QvKnYcY7S8M+/QWTWZHSim6qbcfrAcH0Xu
b20pJlLsZDdjJ6MDJ2oOAqXp/b2Ir09kDqKz5k+m1xrnvYQbPLREhSk6LVnYBr1V
HK/zEyuEAfm93P+V67VF9G8pFFOG/BBXJYboJP1nCEwvRirIjtC5nmp42UCE0RmZ
mU51BeQpdnWv2bvNmuqUtEj0yJ9+AgzF0aCfNBAM8otedxZyEFRsbMFFnUG+4VpH
BNns+Llt+ZRDr+Mr5oTqUCUiwSTa/Ap6dxuWxxbMQF3gFP4IQxoRkj1JufbWpsPf
0EUp2IjzUAa24w0sIeG/vGn0JpYTfn9ZTvftyUapcyMTrF6GHSGXNr4TLnOgzXg6
vZDy9Nc8lvNgYivIC3vjvowPJkyIDLyUuHJP/8FTO72bbz8uVdCfY2A9Z7PFHSiS
MAgCe14s5pUfd/PK9FTT+u4+qUx0X9t0xAeuzSGEz15MYVvbbka8tF3+emtxlL++
vz5SwAn9M4yCglVukVYBU4K9Il5x5DSZ/tllMS8V6DzHmf0xh7TMBHzfcveVutQz
4et98DUhOMjRVlPCBJjaW1q4C+6s1CBoHvzoNnWq4HnaFLY6lqlvQXfnGB0b6ahe
C+U8ikHsbps/31LBnZ5OJ0m+vuPFrlBaR5BUzvg/tSEbhQReQBYXH/4sQB47GFpV
8Yi0JowmYvMgEZ4MIK7CmBrNzs2Swo8tI/Nz0ervZ/XR1o0KHdKoW5fCjSJevUiK
osuz1xkWKUwKbIabtrWZvvPch+QAXOY2TrCSxA63F2kNyqCmUvMf/gQ/G/tz9Y8w
HI660olrXku3ik3wHUJpVZCmY3vqWh5GAArzBakUXSI53zCODY5UUUdqxR9oFc2v
NI5Cn/NEmkz3UBo5P+z+Dw/Ga9NISPJ4IN043BypKfKHUFXvVPSgCY2FFBrpFk2e
FgTBmV4OjBRKQl0nyb1lTfK3m65D/T8muZfr+Vq6BdqUOM/9coyIVXFk00NLiosj
ss7nLd3D86qVCwQpFG34+aiAmE5+cel3HYuVFPQOjP7donqoI9ojOh1rUPmY7Kyl
robtQtLEtzjRIDmf8m3n/8E4lHkMedMz6FC/Pa1MrFzEC8yYBJQDZDlZyXqRJd2V
VZOY1TMiUpEnZPsIqKhe8s/SyqHkh5a/unWRyEgjM95bj59764UgcnuUil/WiXv9
XGR6WGVySSiNF3xo4v1SYJTz0uugwEhJh8dtVZttPeQLeDV/dCJ2LKbeA5TJA6xx
ivJ5fRHVnGi6ypWJ0IY9DbUHx1QS+EgkQzIQYAwG8J3u6oY2o8SucZkB2JjDB+Fe
/T+npyS0vYe269+jDqeWhpnJQhaTF7odixOKDcbhw0CIfOZSLlK2H+qdKcpwCxYz
1u7N53jdd5KQuc8yxEm2nqzW1v94QFB4gWaBHlMC41CPvncyBBmaGlpgnntdYUc4
8nAIdD46sJsFILHxPKZ79h/y0uKtSfWPSd7Wc3Cql+l0SS1zK1Q4v1l7cfNLvjRk
/hCzdLZe+7vQeHrmu0qOZoEetVQx56u5G6qFeCOYKKuoNzLraPcROFcrb8ososw+
4YhC1q++EYiYeZZAwWJrwyHwgc5xBbLap9+0CAU19/1M/9uL5EutaPrvoOn3DFFA
rggINviG+WvUgpQ43IdjwWabNq07LFjYxf+79yr7o/h0mcM69Zlk1V1vJQ9cXU2N
/y+jRUQcGwCa+hkchNiUu1j2VzLC+dl5POyWUY5c6jcuYOufNsq8J6n+CKaVUyHj
vRm+8FHj04dRtdR8jWw2E6MY1OIDRdn3LnHI5NAzN936BTyCEpNCyTFL9QUSL9QC
drexGA6CBp5gib3oEXh9n3Ajb12J0wnJR4KYggYMsztPXFFbcRKfQjJMrfphV0Ad
JcQ8IC6piHUZwd8cASyCba14utWiWfrt0OwDgVsFkkScvc87dZEVsddQucvScKyV
i6XcEVbq8JPs2ORVqXhipcnYQu1jec7mQ9utML8J9TyXYgYA+3czTV3AJyQszvox
P9AToMRf/tVgN5lpSzeBX6w1mTy//eTBHZB528NZFoK7lDrz5XwFBWlHHX30/kto
ZsSYsznK7s9KDLvu6PSyHJcJ9+v+sNNEERBiwB8Dekflpyk3j1ewYv0tvu7WU8mu
aQ6knzRp4z/XVlQjacmSOijMUUaFju5zD9OCLeTOYGzF19CnWQRzscT+3vfeSzTI
3bXRBm7koGGuCdcP9SbZkqgeJLaO1g9bqcKWeHhKR+cHCJ7Pf3+C/iqbanARZZzB
/6tkakAzM3sS7nfcrboTLB/q8vuDPWlPGcgQWEK5dPntL8Ut0SA7GEbnKqRCgR7c
L+HQPL0ER94ynkbCd+5wc47QP2gH30AOjNFRt4APQuHqsXtvLfOX+nSPpYlOUgpK
c2ok3M5mFDzIwZl2CU4wqaJpDUfrHhM7/alQGCQqO+19q3EEdBZ+k/jhP3aLAhcq
3FS5wUvqTXRotTX3Fj6bAPvsw1zERDFYIr1N+MmXNthM7BotgdcStD9ScknRU1UX
IOFAnxjc+JLs2EMzF45M1BBOgmBvNA9DbUH3WqexRT3Q5V82uwgloojFParpPX6O
+8EmSMozA5a/+cLG/CT1iMPybwLAlHQPOSRe15KvrO9ljjqlvRzayyI+4GV0HkkE
phLx9QiL2/DDaQnv4JW8Eq4ejhawuVUO6Qn5zk9Csnknz9++GxNmIzLZDhe6iSQ3
PZKUcUuFcxq2sy2hMPlgIjRPgOFqtbzbO7a8mQETpmdmZe8sQpYQHO1xZconc4vN
3+1H2YMpWjwlbYK1fAAFX+xcusIEGtlWbIxnoKwtN5ucKb9t5QvVpZ3l2DlRZ64L
C9TSomsYNxV8rP8UvY4i2ZXNCAkCDtGR18+qTCNVb057IZE1tSjs6h9wacgYSQd1
NGjJ3r6AnGCyGmd3y/aeODhI/2iNTQOtDvKXL34KIAp9XPmr+NVPBJhvKj0gk8a7
D9TUhlY7KuciO1rrvXRUglkUcG57yRfszgt6yZn7T+ior3moS7R6u+u7MDT8Lgl/
ocXO3Y5cNvarGlG+UwKeUFpSmM+zLavX2jfNKI7bTHeju29SyfEragOS4IkU5PgM
7PBhhLJeyny86JeseZFpZr0Vz1A4Jic2L3ZRkZvtYkJH+GsbauKgIWOZ/66TszvB
j4nCIIDCWhmFGLQFRZJk3rlLfrTp+aqCVlCINyYl4wphNCbuhpnr7HUjerVt1fDz
Bx76n6ALOK+r9EMCOwMFLiaWVJq/jJk/MkdgOKrkTr52tsqUiL3p3aUgGB6Esa5/
UMA5qeWzdoDfDLBLeSLaA/vvwvy3NtJJgBbIr5FO3jkSb5VsPTKt4LK92FPMLq6w
fkVtH/KjLVq+jy8bjXqidP/5IdjmQcYsBZ1VEIpPQ3AteLPRjrISDra2EztzlLBC
iQZKFWtAJhYbAcucQuPeB0GdkdQPHVHAAjuP/9e4en/DjqKWGKhgpIx9WC/Pdrf5
d9TzJR1gtcON5gLeVP/Bwr+TBIl5JmTzFgP40qW7jWZdydS7jwzN3aFfORy82VcW
dXCNrjgCddRmXS1TOuteRXCXt7XeLiLCfM9PWANHb8br4n393E18ithgdWCJwXDI
vk+jrleJNfaadzn7gpiLb2jG96kSw3l4NlFENcp+uBH+xcavmkKsmyNMYxD4d3S9
yQZ2N8CS/LA5V5K2UHjp2H9bMiBlhNukW96RnD7LmXP37whKo0Ti4uux/KW+6RyI
EAOuL8UoN0ZF8xsDYK5YPX8YGnTyfrIuGrMwTtKx7wpvvr1hvUE9rrzcGdweiG+E
nheP9YF0P5QkBNOVCCA7+4XKoyj38Cj9T/QRDk1XNfgzcGEuTeiDz9GO0+Tj66eZ
+ZG/T50wxM+fgIRXOWq0WtfpYRtrVhMm4stGWbvaC1sw7oOcO+WG1QtLrqU3F8+z
xpmMyiAnLuiOMFv66teWiEImkzoiHgFukhDrXdtjE5MipxoGsDCvH3iprmgKsieI
V61JbuH/9w9UmjaXjO1+64DJ7s+GoO1GeqMZevYAzuwImRktU3wXrNltfuzm10Ik
uWfmVmBhFw1VWNDkJETcQtmvxDK1n1pSYYEtRvqHqV5RMdvEBZDNof9evAOG8C8F
bNxpQZVGKQVeJlRb8L1uks4EqUjkNlvdtqOYSkNAe/Y4ZImN8/etpk8UMddb7rsu
25tK6/fxcMwzwNNEr6E3g2HVz86D/8utWs70G9T23SmzGtqG3kU6tl/zJgX9UZE3
E9hvFcGMxMGwTEbg7H0lT2ly9pbx3GZh/1TlcmIlXffxwFXsCGKW0XwMo6hteBb3
9IKrk5jeXFLTy+1wnPHfWAMIlKOR5wPtZFwva8fXF4VxhlLPUJ+y51tMIbHuCTR9
p7DNfFUdo01yOPvvjpIKknc6ESxKXF2msxBjKxlEk6libBEfoau638hH93d6UhXp
2YbF9GjAAgkH4o6lD29EUbUrViHAuk1Ch/4TgXqHQVscNPw8z051FOTqAJxqpwde
g4N4/xXPm/erriG+L/7GPe9aODlNfLJyhg6+H/zCWXwtDxlv+F7d4rQtLkfdVvIW
lAHHt6diZBxMHvdk2Bx5p8pSDzIYqsnnrJnHKaNqsKdxt2tyBHS6KICJv65HCZGA
ORt6kF6DEpHsLzN8WItgFNCuKOjuKP9Wje5D0q0UCZB7NkttbEn47tjqjZ4Ohhcq
5Tj0jpnxEgGlUHQEJntk2bIFMAN1aCFsPqtLJXNpcVvm6LIQem0Ccf3Nr+8y9QpK
zxy91nqrILs9lDBjrA9XE4JzTrpa8IzegHwflnHmgGj1jdIb2JdPqgzPk2NLU4MK
53uzCw4O7rRU2VRROozGAd+e47t8VLo7vmwSHtJ/iv/4tcjJ3SpFP27z4Tux8Uvg
ETh730BMMBKA0gCG9ceunpuRsD1v3JNTo1ILSCg75vXybn3o4QTBKZFrmyg+V0NE
svZSzzN/kcQtJKrdpB4+D2drtXH0CuI+SN2mihsPpJncXQm1e77Z1f47D/tvS2VH
2cE0PF1FmAv2HBxG+UnAKwjzBTbhqWmi0gbd+Q0P9TNRwSegL9N1DLIokefI6zw2
E7XX00uTfTJgyuEfkOFaYP+JH/xgfX/1VieD1vSTEuA/1k2sGjTP2EAWSmgFW8U5
sTx+gsH4VIl//eH29lRwcQ3eeNWLpJ9/ztph7Sce8/sRVp4oG+3O5IOQ1PFEWqiz
bQ5i4zS5ueuj1XfXawx7Af3B3V6HwwJf3GBHKxHCuzA659B+9SV0RjME98jUlsG8
0ydKfHGtG/M7Vb/kqtLdOw+1CdKaDmQ0VdmkDEX1fV7N6OlWHIxOH2RZfxomwjlu
rvwrpm8DThwQKT5zxLzOVHwLiS5yfTtLD5vWhL95F+xpMo437kH+3hGgNJ+qA0Am
cePsfeQKbUxrD2fzIxI0GsItzKxZrO5wocjfMhTjo+MPIaujikS7Vm5CjE+DB3lD
341vhYqVe9ZW3eEGJnCgLCxWbfhNpf3QaYAYwPv+ISaBJD8EgS8v/jH5KuFSfotZ
BrMd/+7jC+icVVtIofvcQgD0a9eyfx+9MVXV72PWLRSQfPtpBb9gNsTyQXgEkkuf
o0C1Lq6LVFhhFWHoLQvIO1unuI54k/EWjIUAPDwTKy6RZpPWF3U7klMIJnJ8/v5n
VVw1+PFJMNh7TbsspkOIsSdk9NuF4zSIdH1PAULwXb7s6OkZ1RW5w8hNS63qHFmw
Ra1lGPithUx6xHJyutUs8VAOHVXxCEt5xEgGH+CRDSbQADzONr6HzhUwwe5GRzji
kDy1IvhlGIEKNRhEobagrPaa//ccwN4EqBKD1RFhlAjv+LC0Gev/j//aR7oygrNJ
Yos+4bvQxWgx7UPu+6KMrFtkiU5V1diK2p3dwQpt1ChM63u2p1XW4xQ150jJ5UM/
VCdpjihxUBy9S3opMGxmGEv3aQIF7nbnL6UjQPeMaVPGO6gX9OFCoOW4WltsWu8M
FJv7iRxQORkvBsloZpTAbI0HAHizDvm7bCrrzs7Orc1pJBko2RQSSuUGiDr73EBg
qSaVuJMmxwDWeplHij6sXuEk6Bx5QMXp5upan9oJs5r7aVLGPNyYFtKvYfikO1pG
aUNVth6FRCTXz8JGS5RvOaSrz1/IGnL2Pq91sLP/6vX1yWM99NH206bHDzoIiiwv
Aqtp0S5LtnBgde04k+gN/426P6mE/gn3qu0ZdnKtlL0KPi6OsxHKSDlhn+ksIlPi
WseC5kFlQhNwCvuDVO3JAJB+5Cv0AGlTuBi34BNDvC3G7ecZoYeWHrW45fN3Nnf8
pZkH+dqjy+4NIzTP8GGP2y2PDBus1BsJfje47KU4nmbgRVpEE/MULyXJqMkfunOJ
V+D9iY9GOWFe9tTTXWqS2P6LG7XDkZ7GXuu8IXrbNeen8UkkWhlHvSyhmP/PTbwI
5Pvgqikm6Ijn73gfqzZbDexwG7FXhCL8Bk3gBuquXWqteFROpl3hmEJMYFZslr9C
3aAQdsyIkBg2FUKChSM+KERilIb1k83ouZxIDvPiXmqvQR1MkSnaM6vPm5l/+Uth
Hd32wGHdqY8Cbb0kbyR2WssQ4eZYs0SaToqeWprGZ2pLozA8tc85MGBbnl6omeQG
tKlnTD7EXY0gD1IJxyA7Pa27WjcR+r3JNrYf20odH4v4E/21bQ16DF2t2/QlWESU
03Z/Jsm4dSoXkui1x8H9l10FqJ1W4CemGATDZ47NPvQj7GihxxPYUQkBT0WMI6mF
L7Yh28W2V8RHbn88scmcd+4wQKBbOLR+KMxDRFXyIPFOJav7TzLgvYIh7hQQzZ81
CgZFliQWcLBSf2HCZlaCifh9+zRohIifp0sSf1TeyOl2tnxMwUmCgeO7OTdlucBd
+P/zrLOV75+OQ/KM9zvTuQOI11QcjUPIq1BgIra1QXIvjWULX2KWrOPyR++pRjVx
d2ZbWMsCNqrHfSY4PeqmJ5wLQlvNRCTI3dsq3dmD9aZT5fQXpm8JHR7AKQpa5aQ2
c930oE/7vseUIMqkTab3NEvdEIpp/QkQPXKT5kB27kAjsK3/9LFH7MomSjhYwFhM
n+ZiyIdnrBtvNz2mZlHdPE4Bz+Wav3ex984z7DW2Xluwtj/T/WAZnB9X7TFmuA2E
CMHMQUA05Hv3h/ae3mCKpPmLbVDl3MbpwB0QjO/5BrD/USyIAqJSgOC390P/kAdS
Rba8lkfg9KXVRaWhm/SdLzKBGkvJHMI72sGyvgdgiLO7F33Phys8blkhppSx6nf6
rFEGtjF0Dhgb5nNyjmhgbUdhOh9Zol4kGvJO65jFe96V2MU7bcq/UDAEzA2lxWng
Cr2dVl312YlN7bHPJRxf1bdPKNgKUhWB9PIcd4ZG3B9A8qitXpAKKmvoSbQisK5R
Y3nc8UgoBr2SbzKFhY1J3Qn9YM0+azxAfL54JfAjE2sBCh0zYlde48LVsxr0Mb6/
0lquqROZqoI6wJx2w5fRfI286Dcl9pP9Yz8jsWr3w1eBtCroFm2JaIOHeIIhFKbK
Rz9pOVwImmDOgE7tA7t/v55fogpmCQLQ3ZyySpAX6Tl3qeEg9lla2b2N9Brbz459
cCXgKqivGPxoOS54D7ZXYq0RF4Zy1kcnaedzExVIkaSYklb+/O0YCsP/k2c45abp
brkKIKA7ZqF7EwPqe875pQ7Q0xmoNVMYZfbZEz8ioMl3/Smu7tNgdXylf/aqECdj
C0U4FG6XTrIID1/UoTMzX9Xr0Kiv8ei6WsCrQA7W2O19EwBGAM0sgHV9HRjuncfI
T0Pgj+LZPCOaEjStZlNoXLAK4ecSjHSf9U2RgvyGEsUONeJGSd3XjoyavgGxXaW0
dzVvUhcoGiiwMtZoc6fgFQCb5BNbrOvnFzxnrti4SID1PMO8aNhoz1xrd0JiTxrZ
xElOeBNq0Hxv0pI3NiUmUInk5jg/btNXZc/h/M7f+Gn5GC8W9XDujWxFfXr4TUo/
3nhmNmJcLaFMAhEAzE0QUpRVW6c0SuTROSyLjuhyWUXKFoVvIq1dyEtvDW4hGs80
lRThWypJFhl6ePtTFgXauD6gGia27nR6yhiVKLg7Mra933D+FmHKzgLTyy+tZ2yg
SyhUWTZccVHimTadnNlQcRYSHTmvWbtgF2pOmMLjpgXLaBGC76MG+EFRAUZDczG8
7ObSve2feidnYCO5lqfzH/jsds7+ixsqpYIdcVYBe3Ai/nIz6uIiz66u06UcowZM
a0VwLCnSwDWK5nhqcQFwyDkwiBEAf+XZO3pHpl4TmaJXYnwy9zgjgC1oVMLausJ+
Wl06m54/Mbyu1ZXMf99Io6jhNKj3R7+fXTKYDiTh/ddLaIM2D7BkQajjcp6TO6qH
g05g32fzSLD+6/NCHIA3R+Dd5HSFvo47nX7YzWNWHY1pS7SW47cMKB8cIN8t4aje
3hSLcKV2LVjPVhs2/GUwbQp3tmV2/v08RJgFT636jrfVf9wNqK5/iHBRUshR73za
2sFJmpBUSO17HczJL1i9kTq5kfDzndhZ8kUqCmYUcncWwOhCrjbNZkpWuopKY9au
qOSV5yEUysbl1ZmRtlNrs5Ntqg0Fp9E0PVwlhiumxDFokhjvNGavvnxHy484W69+
mmHM/DWGGQ3B4hEE4w+v38xY0FihUuiNjlMRtCWYYuRd1tHUzzQQi/XHMcHRbr5O
iTTuZHOhV2pOeW24gf9gy5mQdHNmD6ypJCa5E0j7Q2N8AsvfajZljKFkwcc7dsZk
t1UJ6At2EjzKiknT+w8RwUDO0OVaQ6Dh8KgiYcY1NXitl+35tr5pIiKZVUNblfr5
A77egklv9IHP7MeH+HM2btxcti3dvGQCmfkIFp6Y0l1gerhgoSFDM8AlwZhWqGIT
DrrJUKiZJdMONBSFEGv1/p9H4XWDNvQIIZf+T02VfieK8O8g4NOKshnxxQaL456V
5kWz7nhUqiEB5J/pMohgUXWvyX/zTGAQij8rGRhUJSVv58CXLn48jhzRMdrr9Ayu
RL4eqERCHaZJIedjs8pbShSNfFEFEGlflqXXMlKM3nu8kipe3HOs3KsGqj7JSYJj
uQHB0C2OKT9b2uYXCxPAUEP4AwtUJO28zzy37m4mTK0it32tJVn//iiyc1lwRTS3
RlTNPTxtpmvTrSBZJcypb2k0SqAFYwMWggLKwvgwles7rw9NFdUrQVsyNKQSodHL
ikDi4GL3x9uO8ziZE5qKtbGRSI3qxJAt3g7JUMbzO1io/ivEOS0uSVo3ZaaNQei/
lOU191ZrNgPIq5Z9TQEao5NmP9wlE4zejUbmn83H1XmYMUF5bmeJWJ27VCQGxYjM
S4w8Vci3oWuSP2FrS6xbfBzkK1bWMpdjXolPgbzvPQNumGLNUESQLTy+iVJie0rR
q6bCmjituo5rU90phXajxcJsXXbp1DcMQM+wl5V32pAKhyXStwFzuManhFfSX4PD
Akxp4qTQuGuDvSxl4S1BY7cfSQZf2frWAmpWA4KU0hha7eH2givCVVMzjA3AOqzZ
+VXAFHtv3+VJzrxn919usrUzlV35AYIZmMPMy6egJAFEw2cbm+LF0ZBkefwVwidy
WyV5GH/Z8AK64CJeYhIUJf56KNY3M0M0ymIPJrTilTLcTb8Kfs+fmTI/Wocju+uj
c2qjl43oyKT8NCufiM3+tEA23xxJJLyrjqSWgWFIA2riUVdZpSBB8IlJWhXKsdf0
TxZRvwImrDihfvjrhefV3PNxD8e/MZWD2bXxifj/nHqDF9sxnuo9R5sVRjFkBZOO
08cpx8LgW/TJmko9I0DMd6LScmHh2+t8Pf6iMCf/X8IhI5Fz1nB9tAEjt8Lh1Lio
ErklXurtr8R5RgJjw+cn/f0VM2FaF+dV6bsQg0GFOAULpyZ/bs9CRKFQkl159Es/
N1ngDnXVmkhJnemkmNgSNqXiqmE1Ci0cDOpKPElVFipwqf5PTRDmJGcaAQibsdlK
yxgTeDeSnozCJHWL2l59YT3+11mBrsMwmZFP65ndk1FiHy9mBztRz2f2dVrKIRWo
50xN1LZzBOxnb2p+/35US2D7Dsub8Mzg6s6pKrKJkyK2mXq4YzYIuUWAsl9xd5K/
dG8mEQtn4WYAyWbCyqPxe/uZv7ZZ9V/v0xsr4X3iG5ySnWX3B28I7MOXbQuQkV/F
oTUGAGYuT5e5tNfTWAtl8j2Xm+tyWMf0UbnnSEpBFrBCwgW6PuO5jk5iINt2Esht
VUcNidpByr3JAkfJ7YY/udBDTLtRStWek5JxiWVqyQ5Cc9eFvtUvrEePRs7S54Cs
gLSAq3u/cM1prCza21ShaSCoz+1KGQCivgxRnbrPjoL8KXHR/ilSpT1cQ4pvpyzU
lo8k3rd0dzGxxDbS19TAxwRxSld1waPFeVBHPNkw9T28Iq/mX6ibokXeXq3l3J4M
hKXJS8L2R+DXwlVmYcnysXQxcVhh5HYKunZ5k3Xre6stGnGNcjCFFoQ+6/+fgfvW
LIcmSeU6fH7A+qLLUCxl7pawduBLyqHGkRuj1r0xmYPykQvYP4reDu+Zi7DEF38m
wcqpdy7iNIAa81r9td9vJVMS2snIvRE/NxeLXvAX98xLurpU3K9hIPoIxm4P4uRw
wI2ss+0uIfUjd9Q3hwInMW0Txb3Y8SvTd5sm4WPjUJbMhV83Uf7xDkjaSLOYhKCU
3eFEMh3PIELPlsh0AzVWYdJzRWeLXCoVCz4M7UKbgi95oRnujf4Tvsnu3Cadf/4V
vXvBf/nqU6ytx9hJuzm10zwBqPsG/tElwdXmXRwvbszBoNGbGEJrnhfZEklndFvU
UK4pf8/dgvUj8ZvGrYOl8gHFIWhZpL0dppxy7ahJ4hKqpcJixIQzD4ilE8/OWp19
XB2uj5ea/v7I6K7v1+rP9GsaOQVOd0sUTD/PVVyimeT0lubPZu1KF6EQLludEny5
b9IK9n2Bn7NNNiz5PMDOBjdFVUU935bOA1QVBuXLnMeTDrH7RQzhYD4smjKGnH+3
ydoqca/Mjckt0GRlOSkWq7IaRAiL3EWFZJMjZ+aZE2OAAXNj8Z5Zc4UknTGsW9gk
6EaGwG8QuAgPCdBC78Dmnl3grZQwmzZlQJUbb0EvBnEc5kB2DD8OFY0yV0Xo8nNh
eQGVJR45SI5db4gO4YP5Y9cGbwvFYb52ank6cEgCl+47Mzfj7wkUcn9EIRBgash2
64CVC80ZueufJaRIKkxXJ366CnoKfbekttSoeX2uYbcOKLIe2wC7wpev6An89UHF
ONBU/+sy7GKgC9dj9gErQ2Mp35aCcY8kQ9oVg7m53UMtkRre/iwJPncEZFUR0tFC
8lVk8JAvpJ4TNxJStmA3MoDGITq1SDVSvvVNwcjWHD0GzUv7FxJP1ChJxQi9sASh
GcrlHC8hCt3ju914TQemewer5XCQjZliGh+IPeLU7PANFfwZbEx0Tj6y8wWioUmP
tFK7hmwt7tsSvKLLxI8i4SZ11GNauYUMw12aVnBfQmPsAXpVnAAhphEknFnECIuB
/oUVwpeXvmSM/yTdBdMtKoDojZf3Y9TpGKowc0CcYNmIi4PdMKuyvuOoARe8p6Oc
QnfrXroX98prrIK05HC779+Kb70UnHEAl2a+YFjYZQQy4xGXfNkLMT//J/HiQqT1
EGxHGnD4IjuQIY4m3ikAceousSbOu7CfeFMkP7QUIf0pf5LD2h+GrFbG9rInAi26
YZAQgN9OBjxz5Or00Z1yHbKTtnJoJyXOHnN6kNH4q6v5cskTLeZEDc5rJJPlasqh
`protect END_PROTECTED
