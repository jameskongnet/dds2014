`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HXOqC6F1yZQkx1p1eIf9sQGuSi0RB6nR/NJb+xXg9SJVx/UMR76AyUIGY1jUvjCx
0kceuma9ogbtrELK7tC/XUWJwRUHQ50GCvNAWOrB+acwAxjWVYRmkXxAW1/IaFfh
u8f9tYSE4q3x4D+Dwx/qU+J68fGOCBU7bQcZgJyQwPrSCArAz1mQ/wFBv5UZlwtX
2nnvLTqkzyxdA/9eNdnjKFarrgnrZolQehm2B36U9DE+WMQn69KUTjT1t6PWwOoj
WGl5LU6e5qOXQ44N4RrcBw5gDG/3dDpk97qpHnL5akWP3v+AmDblnI28unINpTBv
pEKfVX9POdWn5Sp85hALDpfqq4pOUjAGe49LpWrzRI4yS6IbPb2wyY1JRYp0f115
tbYmZcgOOzTCTCqivdiEle2nr2GGBUkTYyXddXQLxxrwKmfRDIXD7QxiP9wrtaMd
sjv2zwBEu49iB7FCyk2WB0sS2MO1++NVefPjK5QWUPN+VnJjE/l8QDjTV1kRObK1
z2tbDwBAa8Lt2J/pRwTIuzu1D0xNncjdQx6wapMR/KplYYTG29wq697tg/FDVFHX
NC5o91VDlLCoLMMIohB43IfVvl9PSD/WFNX/RfSU8m/588ohQ6q2vCXWAu/sDR+z
l4wF3X2f8iM9n37AWYIhNc52PKS0XQ7nJj3Aje0r9rP1Rjp6pU2SQJUV0JTGerJ1
r7/a+L1w1fQbrjvXfRJP7NjEQoKh32OZyHk6QX/2UmfRQuyiHWQ9RmoDnOByCpi0
Ywk+JylUW3coFtucaWNnzpG0DHCbzUjWUzwiVfwD8xJsbmGVyBhaDzxRuD77E7Dd
ZIcPqeCv8WMIlbbhTSzZ//AcZ4h125z6Q9ZGozSBt3cJq+d8zXH6tBDUWNBdiQ8+
0wmlXE2Hr26Icqt56npgumuVf1uVOqV1t62U5LE/IWHa2kteau6YVJnFOxf7HjVm
2ErajiaIS4cU/ycOznHsSBgCn1vg0Colz5xmPAe2/up5i8CwCOl4uQSeQ2t+1EYv
uUbTqMCg+J7D9Ja7Mx9K7VC3d6aWF7EnVthKYaTPXlmrox5GxzwmdBN1v95IrFKO
JgreTQLrmCivR/QwwqJgxmeDcUxT+ar8j4vuJPCQEePlTeQ6V+6wnaUX0bYZSSMi
QoYu8nS8zCw9LGvSqZSSXi/An9TReQLlVVKhQj373QfyHNar/qL/wUQFNWu8Z4Er
fTEr6IUC3eGE9qvAGmnhI0WDyQgq+0SYEBPzhEFrlOg3eceKRduF0zP1Hm9mMRcB
Rb60SEzgN4j/NBEaFj//2bAFeQ2AVVCKgB1jEUoK/Mj1N8aox3ctK3UFGNdoXW/w
M6HTQdvtPHjt4VwzOgJ5Q6EdWSAltQe+FDYNatReeZQCw0DJaTvWRJQ3kVv0JHIX
IIqM3QDoKCMAi2HOcrkQ2itxhmfkS60TypujDci0rCwGhF8kvHh8BCn/4DosXfXo
grrG4y0pXS9B686G7mFOdK+Yp8T8HujYbWa5C3ep9D7/ycQkkpyiuXfc2Ke5LCyb
qRcnPW5jkxDBc8RwPGsGtqdMjot3wOkJJ81gjQIxwIUqWA2rQJMBntJeeN560lr8
1O9WQvmkPQVSlCgiRyPKAMoHJi7j180fqHXlsJrdhIEXI/vQpERThgnZvqjB7YHF
ycO1swH9ke1r5cE6Hs1SD166XnYeZyaUbSZRaPfgMNOKmr3dH2hfKCDlFmcKfXYG
57uOa05tJ48pPdW+QeX08V9QTX/S2sTLumNYDIo078kiiaYxVYbU4pRKVuQPrQll
xxokI2OfTNIU9A6rFQkr0BO11e+F01wPazui4DNvaLMEjD13z7Xvm7wKQbfsIlQJ
LRRXNwU3hJ+zuCNXu80JpEdMv/L4qi8IWqy3iAJL6mWYXe2mfgnM/sMVBJteGhxy
ZEKcvhsDF3tXcp5hldHf4QmjXaiZhgjBNAfNTAhheav6PnXZ0hr9Ff7GgZpvYPxD
k6UW+XC4xRu884lSZVeCFt/AUTEwixtVSRxXYGP77TsN0QLT9otWLehMvYftenkS
GRnA+Ve+UHSJvWlZXyP3n86jhsb/3fmCqf98XEZ3Cc5JjF2c3UYcSX0uZyrLMZ02
d5sYjNR9M0/fbuiAIThP7+c17+lxz5LmwVe9QHAdtU5iRbDTICmKYpS8rny9TjY7
7Bnko+R62wDo466Gb0ueB3BqSTAXp60Kcoq294RgpBETwH3ouF9MXcS4vmOkKzl5
B/DlSQUoJoa3DzMu0a84fUxyDRpCng13sBtnMgGxgMSXvWYRW5MC1rLt2QO4V5vI
6PHTqMHm4Nka4M/Yuf9qU9f5Sw/53nLSX/FaYvKwxzC1UnQh7f4ivzlOczXliefV
jWCCQYVU3jd25eKRKMoHNYcULFgr7xpUU2wyD2BzTjerkl1VoEYT4Crqdhrx+KUB
ApsJl3sw5P2Pw8p0mXJuzYew9F/3eWBlBKY1XWfY9w4Yo2KisbvvjhqO8IbY2Mri
BCjfDNPBmkG7vdcqz3jCg2PEK0v6qVTj/o7tWY/46xRmDEfwaDqAjmUXFg8btnSY
45vEg1cIwTXXEnDMZOJiVnnInF8lol0mMJupau5WwAbEysy60LTTBc56N0wdHFnO
KrI9WKO+OeFOK20DsoY/5uyyIUfu1lrUrWa+xOBJcw5VaTiTzL4s3eL8S6O0dUMr
ZHZ6794Egw+ZUUZeVNfGvS3kuuRAq4ZCCFOM84mg0KuW5XFvt9vEI5+qcUjwvfNx
a36EV71sIWopYKQm9kV/9I0hxGIXcXERvP53QXKb0ILA9slDYTfiCPrNTHcbhwiT
bunErq6s0q8CyGE1ENs7DpOAly+chNA3dt77TwBjX4VwxqBFHxRWkF+W38NPl2lr
uvXyjjSguL6DRTIoG0K9ar8uOCCH6ypp9zEsGKmXU59FvIiwFgbqvm3Ww+QrVEAd
FipCT3hXM4WraNJKwVRDc9bxMR/YLHTbDXE6Ltmj531hmaleAgJr4Qn/Bxce8anb
4tHLNnEpZboEVILOlXgN8M7vJJAj/DNWofYzWuvVNwwDn0KZsbaVjk1M4WKk6+M3
9wazt295J9ufmxah3WxNcLDh5+I2mYIVDMLgqa8xWGXeM1JznjnNK5AhsO7fhdk8
UEd1bqk8pYAllki5OfmWjB0/B3wvjWC8AOGf8odFrLcyAtbh9AxYveQJCl2BY8Bj
S3gWgxEuQhWxxAyrl5mXRrKoKAjnlvwemZffKwQq2ISPGrOWb/azqg8MpK67Jq8S
HEUbH1K7h/xx87EW2DvZfXGvN6tduRI/VV1U8u744JywWNvF14CzoMfmLczXwfPT
murNuYlle5sWpMSlJrYD8A==
`protect END_PROTECTED
