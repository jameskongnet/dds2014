`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ysXIRAohmQq5dGdcJRCmzMBP1Rg3cXb6QG/J6G5qeWzfpFzRLVnPq/GzXoUdj9l
/N47sMwWyhDvlGg0s0KPJqJFXUX3t3hs43TWlkLQi+OWLtlCZAXtvCGHgVI5oYEq
+OsPhsGoLFOXTZeloNByqUYhRLDh7loCLa+8cjoljXmGuCXH5Fa+b7cAThxsRBmp
53mruo7VAX43uo1CumFeWQfPdY9dFGz326C12cOelLYRnaXVLMl16VpUrbAZsoE8
VVhnlq6tlw0NHb8DTvVoYBlgEy5gozgsNqlNe8KH+AFWYkTDSmKFSB5+hJE/va2V
7R8oGrdWKlYhwkL4fZvDTuCE7it5WabT6mgs0CrnMoxkZWFetNLFfFLa0nXvvMnq
/1ExWYBdki1SMbeAZ0jtTQqJbtA/2n9A8MeZVGG6pC+875N7dISyeSZO9rCR0Ahz
8V+XuKTvaxrxc9Z06QYDw1IVNT3kXwxJP6RioX964Zg+KbiyTZxHe+z/gqzNCtIc
iBGLxrWMtsgMQl06SMTRA4fDXa1xaWYUIJisyZ3WI7fcgBLBhrEntgOyE3BKN+5e
50FqTM4yCcGf0rWD+s+10laF/ChgzRLnI5SXnyIWPQzd191EXh4XAk08yzAmFwpT
cVTszGKOdyKcDqvnNTRT7jP7fk+Veq/JxL17KIU+DU6ZOH1qPfcmaupmj+XpVtHp
+qugIPIhern05yPmW8r+UFOdWix7ZRaKSDiIQmJkU4u/gyrWySGm7AHxW5yebMFL
fWLcGyFW5jPEmFptjTg0UnC+qP+N2P1ulgPzw7xHki/I/b+gZmOjJl3KzPBFOO/9
da+BBlifw+/uZIL0NFZNpYubfM2GLrPPrUoHmMAs2XqYHnqq63BmRa59hizlqmHm
5XYxa9kjd1sHL5AoPu14Z4D7ShenMoGuXTQl/X+PVZNnpI2tyd9hCaeGzVDqlhaP
61yt4SUh1/CpvBy+r1yYP7BT0JT7o0IAGXn2IUYAxqZ3Lv9q5nSbV4i737bxlSv4
AurG6C3HF349IgY8iF78/fIgmTXrwCgRIWft8l8Jy/0kAqhX9hPXwpFPx+fqYwPg
fFt5wEvK3uKwpLDPW+KFofJxasuLYXoyjA3tQ3j1JZg+hh3JhrAzDeNSTlzQMySJ
Lz/7DQQp747QswgFLDzUvMJhFUKS5flp2iBeKvTDstEGvbjgojZph7xMTre1nXBX
aBsahAQiP56nZY4oMzmgbXdMYCWO9VqvkN4wQDA/hgEkfHvG8YdaSF7zcAEW8T3m
GMoyIRc84P4YW8Hq4Z4aGwNBEWLCIb/Fq1HtnBvHO+vGQ6L24rb2xfCxBnX437QW
V7kS1b8zjRbbIjQ0fqpO8iuI3NKiQlyKdoJex+ikegfRT2wN0B7R6+45saYm/Cz1
NydBiBnbWiEj+uwiv79r1ZlGlnoJzHOio4xSAEPePcb27RXNiz/N0VXIrzcUGw30
JCyNY4QGdsJFkQYqi/YrwGFbauQcm87aBHZV9hKgcmMfC2fkE1lHWNpjuGLd0+14
CsqEU5aDJNSmnWnEyPy6UV47wUWY3iJhtuyivGRs+8Ot0ke2D711ADfkDRA/nqmz
7c4dQgRdBUzdCx/qJs+SVyJ6PpB6ugo5HYuaJHyIbw7TxRaJVx6TchcyPzHLPc3/
TBnShbaYtNn2lKnzJiK601IXkWBGS2Vmx7KWVTG/Pblt2XpFBO4+zLMrXb2xLWVg
WpaTSNO7oS3mK+jqQFil6xWnwqiJ2dlopbV+3t5rl7t0uFn7KhUQqYRN7jlCS8EY
eZdhpvuTkYNUjaUI4d4d4qTNt/od2NAx81wdK8zEit3LXpQ9DyH8E04DNWFvwAfQ
ik2JpupSqKb6FJethop5JGd+myT/4TOHb2hBpUQZTO4+Vseelt/OsrGvfOOyQvaa
vJjN5v9L4fzoblyDkNBEc1n9B8WK3b6NVcSEn1etCDMRwQyfAAWksH8UVNTX4ZGM
Jw5GO3HCvmB3Cfrh2HOFSIT97VL9NbLjfr7n/ia66E+qy70bkqhoRPmLrJ0n775o
uXpIApKbUnsxDSzqWpXZUpAMwlMEEnsnA5cV6Xf7PnNXIIUkwrrfK+m+dGMj/7r1
b8Vlwr25sG28mlQCiBawjr0DNLcgHUgHLCfoYNzK/sflyz86u7LM+Z6wnl0mT8Xa
8yQCJXftBqwkdbXoEUHPtILtWcvrKecXiYKSIr1SSOUl6z6JS0aigUCCJl8i2PTL
7UbmjbLNWv+LMBchf3CRIj0fwuMUnzFnqek34ZTCgQbI9T/gTV3UZAE2wHHik5Ih
pMC9QCA6icvbGn861WnVBGqf8kfFknqRlwF5gnYlzronGa0q++Q301jV69O+42rT
56XlB+unroKdnr067IKY9lpcAF2RWSGv79VhDGIMSOfXbcx5BEmPZfK2TUyqCLn2
eGbWfNM6qLzkzTGyRKuIfe4UWMHwfWIXd1C6X/i+gRusGC2yb147E9ITfK/JZeYD
jYNZfkUgwznWAjTeuXrDMd6NA/bYYhwgpEWcmHXBeqUjJy2/stLHHBKbECieGimU
lNQBeBZAlQzt4W6YKhsmeBwwG/wj830uCHu3ONWX4uAKGTA3XxtHC1A36DO3Uvpe
SRLnV2WbUEdqKeAdUcWp+6YsBtte+mbfCR/xL2REhFGZHpTJp629rBQKzWnzFjRd
MayJQKZpoWPiiqPzs+rfTvU/0ELVlQrFgZoZV387TuxmLbY8mJMThc8UTVZXQ/6O
h3JXI2dq2C4omrpxvmtvBBL5SCt6PhzHFBV+0Uy+ajG+u9bZpYF17U1A3czErcWk
rN4weB0RANnZVYaObo9D28J2bwrg6K/nmsnas9DUB76Kpe9Z1ahhUBdsmNSi3WWE
tg3koMsvhbvOkXYvRMuSCWWPAoj50Mh8yg3a9DdRqOdswnCfcnM7Aw3G1T6euQc8
UT/2ejMpkU/2KHwleCtdkdspSAsehBOqsiEl+dJuo1u5zR0dZKq3vYru/BjxA0Ql
62XGFHFyoVSpNuttQSQSoQ0yzvrR3fXJxaWjSE1TNkU2I51KnK6J8ZtDqeuS3F1R
DRGW0bBehKvlQS2MRA0+o69u+2VDbIVXWYFf//vZjw6nz5b0gU1t0NEeco6ykUpg
IUySanu2nuYdIx6ybghuG8j2vROhChFdJws8lcLCWcJVuKy54IqF/CiWFqzQD4/Y
/V8N1yAYcHHmuu+gYI68Ie4KksQMptJcR/+cKQix5E/Vepm/gVKBwIv+/PdFLhfx
lKjuLFjWbZmwv0fzq19LfyDyoGmGhNqFbLRuy0M28lcM83GSAjMvFtKjIRF/Xp7T
GD2s+UAfjqWiRWNGIuK9R2qF0XR26PLolkUWjF9YKaoCbmQTMbi2RFW0uu10gmKu
IzLQe4RD27LEAzrcnsBQF+mWEtC+5DfBdaOhyBsTSIt4jjARLs+AmxKF/uTXc4vR
vEY1i7jNB3XYM2EQBIvUXQP5bSSm9jGeGdR2A35PcPpKc9IWC/R4HkIrqA1A87pj
8wrsNNdSEsambaFdlGt0jkTl179xcBjJ+F8gP4t9cYgjcThEOv57Dcqa9xuBta4+
PXYpQo0u/E111zN/YioRERLFnWVx5XSscTPQl1ThVnDAOrYI+/WRR/n6QMdkO8oi
Zl9s795E15Mc92mztuisbbNrrDmqokpRzSUbsqZDYI1kXi9kE+OT9z/YzNVG/fQX
MskUt/jtsPxITf5hVkuoacQFfi9KYbQlTZOmRjk07hVQ7f00wIC0QBIUafluF3fu
DZ3znkki2rr223q+xsEFUf52eT88s6dEtY08GQN9+9zUFPXJV1OssLpqOcyON/kt
b1SuKviX81x+9L2x0/6Dvi8JrJyZW0dUMQcK8rAisLsqD5lEDP+9DTAx9ExikPmZ
`protect END_PROTECTED
