`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W8pVNPkLETn9UCrQVK4sZS14BmesZpBIY6LuWSTHkdHmkG2CA39lcFz4Vhep/60C
8CJYPyK+POIR/12CEwe049mbml5N6Fc5tAlm92LQ24mWTSkYzHZCpH5jdyApN3Tb
y+goXnmMmJdWulg0/VVIOvykSrmFbWAJIN5jwprZFJVYnd/gaFZ8AtwuvoB+6B+C
eRhNpOEisA1xhcmeHbI+VtFqgxrCpGR6DWgWDVMvY23kcVZzlBwkuJfVC6hCrwJT
cb1W3yhxxHQzvFG9o+J1QBPCnZVMyLRarODZYvIKhEqblPYKIGe99SMe6E60Y3Ae
YInHDbNL8BylfOQcLSIKc/Dq6cAi3d6BwJKKSI+XCNEnskvYNlehi8hCHzTxDv66
CHoyLQjoyir8JV7i6LG2rfHHF/2kLgRJ70STL141rz1YRRrpuImxi0FJ0pfPN3mk
SOm4hmwV98QJGMpDTZ6kVPn/Z2Scov4BIwvIcxbVzgZm6+3R4FUfBeDTvl1o00bd
fSZWmhvuRmRbcsEzwirW1E6vU9sxFR0lLJib39+LH39eommf7M5kzqpMfUZk2Iqk
ZflKjC4LsLBimOgNH+WlkHi8CZ6jSy2V4ptPz3BViZ+t1ZE6IfY55vW9lTuV0c+O
CWmkzTozKNGH8J1Sps1Arv6wkoXnxUWJ7NiNx9PZHtu3rt47lc4tcbdPHGWS2UMe
cz2KTqbW5cgUeCE8Ea538SRQL8Fv195p7DjkUtsaTlSXiJb48rGzIqoWkbnn9j2b
ato10pOJcTOhleJkF9QkZl1WnWRRd7thE1Dxr2Pnu6YDlLEW7AqkT/MyJCYSSeWz
aCh4BObPCNtjm1ZWI58uc+h/3TLgLWguco/4LdD3YJ0RbfAoy3rGwPHcw+qoX4SJ
ddNGH4cD/aGkIxACXf59CioxGDfF+7P59BGGxYV/lkqHdirSlWFc/aHlyQPChi6c
1EmYfzk/3KO8ki8E3SpFe+HPWA/rhcdB1QjO4DLKT4h5yBjlR7Wswmw6vobf3Rh5
rFZ2P9py38LOzQvHHjBQzoSvwU3nm0n0HUvi+WgIEMVnvcrYTqIjRoGgHeo8FExS
3AdeocWEm9CJNWrOnFJO9A==
`protect END_PROTECTED
