`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SLN+FKzTGoAkAbEqQ4ZiUHuLRnyXal7FuSrF3B2JJbX3f/mB3hv5lQnbe+WNCNcA
v+hfWdft8+yCds2lse7D2047OYHVy2UJKDtt7ObquEt4bwbhPaz6O2cWiap9bL6P
W3hVJv+XMs/oP7T14fMu4smXuIAy75jirqzZbHLz7g1KS/+NmINfdMEXdppZaFCJ
i+MF0Sx7+Ljy7cSJM6zOzLAM/N4/vV/hTAQyFXxxjmIuRvY+s2sPTeBdI5TtFoQ6
vHuW/hkKLr99+KrHh34b0xZ+B6PTrCkwWSY8RbEFGkEJu7pp3cM/4jz7PUnmD3pT
ovI9n4bVQvIe5s9uaNxJCqWQWS45Qcbyy4vLhV7CWz2VA9fsB4QTXJbjEdP32kwf
DKTqCUaG7/vwy4Q0+Qlaw/xReZIdGFgGei0P3j5Hf0X/p960ds16WlDsmc6Auz41
VH8aoyTbI3gNeDpja7z+zgYH1R4wqU9RhMmSdEmdEvqpjRghKfAY/g0rkRGi0uvT
bZBJuAcK3fOOixEyvOxwOQRUcOmwn2Ipip7oPQasMdpVvTh1Z502GlrenRMRhW1v
FmsyTh1cvTCUjZCjvC02XtIU7fHuo6wqi/y+yaGkz+roLDYNJtmU6M94JdGfiBwy
ktVSoJmpNS/sJbmOdC/ZWfn4lJ+Hrp9KcSZBL5IbfByb4xsEea8d/AKcI9+Xp9do
YI08Dua3ARtl6N1arp27WiIk3Cm5jJifwCXrR6B+/ssW/LGC7wf6jmQYdTn8kpa+
8gDgE18B5obbkI4bzZaBKydwBkVC658mLJYArV3SmQZWAqTqVrlYf0nSKoaJup74
dGEQYwBTNOGVKrQnseOlpoNGt21xNt9ZBRKYyuR9xxn7cATXrJ5eDtkbh4oLbvc7
8tJTt5MYkkR+Q5j8XSgckg+bx0ag0X+tJqh2T5c7n/vaAV3a8i8wGLHyeliDijE/
YEDP0Kcb1nPM154ycwuEN2EkvhBu7eZXHbxmKcaATR+4pLJmYWQNZIE0IH6exWk4
LTmdxbckf2elOUAan+8ji+8lS0MYoK4SvJbLKX5iwhtqTIW7o1jlvKThs8lR+8aT
FtBd/7LqsJ7BOxK6jSshfNGbvD/1c+wKJ9UTMWWxgyHzhCthIyX2j47tw3ZDuUCK
1oYRfpr17tbwZsL+L8ZGvhcRjpUrYTOIy7yOf96mGWQ5cYcMj+iA49EQjgzVMNTJ
fnXIiUcsJIYyCkdrdJm2geWw5iRzfQmGEQxRy/ODemUnWkumcRVQM7miowGLq2Ih
w8SqdROL+YsAzmgcs4s8aZ565/j/rfK+Pz+aN6RZIMQ852JEPavh/YBtlpAIfYXG
yCCRN/RuonsMcjz9gv7U5VM4zD+sRCzMXVJrSgGXDrfN+b/hBhNa6H+6ijDiY+hM
257MOyVY4cb4eHbR4fAk2er4ugkOFDnXUGh3bvR71FpnapIM4/A/7yrTbfXYVqVY
3/QfmWlSbak9zKdRvWYNoqJ7wKMuPIJMUzivZL3XRqWnSa7CdJBQX0L6upxBYfcL
yLCkvjPaWEgkhQTpHj4Iuio5Zh0Wv1Ahon4E5lT0wNBcj9Glv7y/xI17wfcB2+EW
Q0JvOYB8AW4IQ+z4plXTgzCOPJLjbIkBxR930tv+0SoZz1Eorj6Rny5FTmOWJba0
mT/AVfmxr4v5cREuPz2BfkpSg6JqgqQvkRQFkGbEtNlf8ndzC1/7HVeSrKfx66He
UBp2Li/ZQstMW/SLm1eMzHavV/AYtQ6pdn4Lf3YjXA9J13RPJVqP0+Zuje/HqpU+
6oCpt4Az+c9lzj3d27XnL3Q+bMnCB9l0QKTc+w9vTvvmUFfhaRHc2/tQiH43LyOY
ZIw6RaD21afU59U9hhHSrQfVMH2I2AgozS7meIMf5jZAsz1qL6Ytimy0OosQcm10
PlKJATwN5QgNm1Ls28bp4HOjQy2nBb3Yw+NbL2jBLZsW94V2GO/3A2rnC1FhpWs7
x5ArT6OslUBzKASiH8ODaXQljWcKeP2nzeceB0OmE8f7+1rr6/GmJO4WUODaCh7g
VOPBdJK7DOje1+fozJNYop3SY8t59ZxjJW7Ye3Y//ccy0TOnZiyB1hOPx6VMT7Kz
qbp7ZEvn75h7nmsE6RhcNq9QQoBeY97lvuoQDCFcVVMMYHMoBtDlHO53jerwdVo3
7YvxvlLRjbSR85Gm1BIvYDbWRzox7H9kwRxMoSwyaliFzA9K/WXNsZfdK7/UGJ2S
gSu2mq3aqKQ+vcxAz+KjWCL6GvEohoLciBQ49W2R7EsWMZ+fAPGLfCoRmtBcEjKx
d5z08bDJIfRPLGjrkheeBxJO2a624cmQjy8NgmsqcOTHNSCnQAcy3BSDlUFn5SA4
Si1pAQCkdiAcEk9mySDeeXwsr0BO7Xnfdz/eDIxRLSS1I6rjKEPLOyLJdI18yHik
EZCnXyySzUBv+V6v78sOfMXnQL2XMEKWjKbhX9/R7fc7HDKHxiQOA6EUImHi0BZc
syItOByXQGFdVuL+SjVhW0VXL8ra6F3e0pbvLY+Xwa/anvwO08Xq8ZsiE2laobTb
C8EZ7sRPJMyMQvQxTmlZNzA9wY/xJXu+RAqCw8tapqDe/kvxrBUR7qd/T5GStphM
kUmbHZ0mr5L73zi7/DJoexyDGzDtX2FcTvNNA/kiG3QoGMl+YzwINSbqmPFTdIjS
fUrnNxBHPDjxh2IiAl7/Ofy/Z3k3nupphEvRPmNk2JfGqoHrdmcsh2yiQippourP
2DEwObShA/WS11zTHGszBvPCs06oedYLamZC4tVUH2R8z8MKJtVrBbMLDV5REyPx
hdGQOGklo94b1FJNESmCrEXVc/yEYQrc3hDDonxx1FnYZkwNvN/mY0dtobfQBRQl
9RzBNGubMHBCSqJp1rbbjT55BkyKs51H/pK2gpH26UJqwK4IVujP5H0p6QQDlInI
h9VSFM8Y1zjZMuoCcT86nxWT8WsRdDEoCyBe6bVRdxHbH6O1cZmEXmMH6dW95PtZ
A5w4PnEVf0CXuLNfce9ALkjIirDk6cRFZHbN7N7J0VpLjUG0w0Z5WgStbd9vPJEu
G1XecVMzh6ygobndURN/2U1x14Y+E79AYq4IUX1oprDZGu0CJCpcJ1afZnyJ++af
hTQ060po9f/1LYMcBbjKA0UikIVrBaLPVI27RRoZ1LWEDqtwPXIIaAKT6KCYRzEU
VKqLIndl3LJRzPktWlofPU43uUeTEHYCEMbrRrMF+5KbIIgu1PdlP3OblqR6RCeB
fGo974hV/ATZDBwU9jCrvk/rwXnPspuJOrpe/ik2iguckkeRhHC2k3zF43ywv9Vx
OechT8RyoDNlSrz5bC5YcQfYjJewK69SGzoc3E8OOCdPrRh+4MenVWnKixUBz2V6
lm2xy5EgVNnNV0R/04HWbAPKRroP3NQP6x2pTK9/W7unbf4oo0pXghGZ9JSO8jsg
oLC/FpNwTpPen5tVJBtZTGInq5EG+wujral+Auk8ofSq/nBTUnkP7ylmaKwSubxY
dnyejAye/XTvNsgHQz0hxYzIHzzxs6ZZMR9UMeRvAldUPpGRBTyxgso25P9XeXq3
3x393qe2GORo1jGz8kDs3C0RkgBtnkLCIv1M3SNhEKCq9DYkvvKhNIc9Ux5AvK2m
ON2avIJgM+wb8WuXEfPf/875dy109H3E7d2NkuVTQTaEZweFoWGcJw/oE1Dd3Njg
9Hr+rlQ+SlWxQphVbOLfTmPucwSYd9DR8M7Hzx7nHeZe363HZkLFWjag1dpnCX/0
biFPwcZo3urhRDVcoCkrGLtsMYqqNx1Qqde+40CBE9pm1kTWMW/WiOH1g19g7CPH
qZnvJnojxlK+5gWHrNF04nlFHN2/iUPHGee2MMWpKc+Fhdq4t8E0lH/yW6BU8F5n
CRKExjaoGU/3bMRE4w6CxNRllXQu69gzHRxAkQj5yu/dTzpBqlpuO7w0oamzQny7
cnmaAfow/0xvgVKQ08SM4A9PERgnokyhUcePwWQXWfK4o0ciwFGaA8BqjCLFn4a2
haoshR0gadSgbE5I1WkWSlZjAG03GPAs4S2PPdEEVTaF3WJf4HcyPxw7ZSqfKL8R
YdcwIrU7xDqTMGek631M/SUbad6o3OIuM+WNkp6eboZtcls5ymnChoAwEEtOhdvu
yZVvvc8ql/x1crrgDgBtHM5DaEWTQcV0IWAbluUtFCC/pCbEEgeYpHWLk55YkAiW
Zi4Zm7Qrlk+qIXiR4FBK16cI7gepqGWrSnjiZDhRNMg03Ey6cb5P2cURbYbUF96m
YntD9rpqrByrXZCyAjqAMwYQfFtOQg5zqNAFB90SfDjg42+xkczkU1d5CIf3uw3q
Oi28r2ChFgCrXaxuk6p2q84POTcponolO+A9sJilwqpF1YxPzJdqhWbgYb9TdRw1
31EtXqbRl98+KMi8qYuG2IoWJfx+G8gixFkslGFlaOE6xSsMSp7OeEMY6NdZLMh0
e4PjM5vWrJMHBKvD9IjBwTwY3ZgpW1k4YymyhyB93XY7TYd5sI0SlBIgpY4SEhtX
+23FErxFJJ79FqOD/XcEwWvTpLpOLRc8pbtjbTrcK7v3cneaxYEqvMLffQul80bu
HWVNPAIhKyFopTEu2cL998AeIha4QnOGGmojcnWDFcIuqqr/m0Kv1+UwJuQf3jUW
7gd3M/fzWysxJ886tPnophOMceg2tZ7d8zUJWsK9jh0BdMKhgK/GbNv8F30i/YTF
zyx0auYuMvqXk092NnqnzjaljR7m2FZXfnuvT0cW7VG3+TGwkQm8Kr8fCwcDr9vT
w4ZjvzHTbiqd50EXYSYXryZQblcAKAAaFkvTJEUZEF2rm6HEkL2gyS7io0wczzZn
8CCICp9G0VYKFcEP2deYa//smRLi/bbwRfQyU+hOStNaFi/vAvML2138uGggBT1J
Q5rwXvn33+BamQjJ796oyg0JXqp44T9X2rq2ToZ1QdVPSePVCkNZhn/jQmQ1BrkK
EBsUAQtl3vYlGdCw9e6zny+xHXM8xAOj3AhR7Q3jw9HjhvZg4hDut052gpHaMqG/
bmrRhEH5SiKL5QYnFMtvyn9/JxIG69GTn6pHHTWpEZEmKfyEfUqLBoe2VzxYewsM
T/IzU4fOt2za6+cZ8yea7ydkF75k7khsc6c5iGS2LG0v5OVAYljCfXfkRGHsE3Ui
bFkxYVxDSqP9BjRQDk5CGEBw40pOJovn8tCAetTWicEtxbF9npIbIj884jAm5UwS
xhJCJCceBLipWt5JRwDkxfxtt5hyrp18nWStx5OVAawWyn4tZeELt6Fcuo1gq729
3IJYRIGT4F9QZv3kEaJm7FekkHsBnJeJzwBaj9wfnZdOoG9rfxGZVIZX1QtxUncr
NPMljeCn0vwsxjBtXaG7yQqWwweQgBWWkb8qdnQa63Bc36UdCeqOPhjNVoefSEzt
qOOmzrjZagAbPfndUkMsFJcyr1qF4yFQMAj9DKtks6+zB9+FIdzznLX/k2UaGCSn
8M4xPbOv51FrnJPKEpO2OCWNswUve6q4k7mRexKsJ936QBYJyyeJNEw6GBHJAup/
YoEYlEK39xsdBsCzTyWMOW67/nf5hXiq5iO7MkIlhdtjuB+hluHnFnJVVa+gpxiY
QZwcEP2M/zMacN8HfMS/wt3g2H8Ab2lJ+DFz2invTazaOgp4hFqR3a8e8bsoRamT
1PYqGGwob0QemdrAEI2AwKwEwAN4GqsNGE9dFtNVsYLphkd4wPRh7QO8Je6CsCuw
z7BoeP4jQ/TIYN1WlYJ/JtlydRoyasglwh5Ds9Qevm/4emwwl2tZYpATt0Y/li7X
J5lbmxHkqIMhBX5WFHaRMORfiz1eQG3AZleeCSW8edff5CAy7X3gb62Z94enIXVu
9/z4pH6V3jamF7iyNSajQmn54nIvBadbB1ldrbO/+rXIMDoLrGiBHKkMJB0y6IAO
D6eZYNORg1eV6Gvz0PXsY5dOqOqJuHl1O75iWx5b3RAgw6KPxMoQwpvGkrj2/PW2
4XbLKBL87h+6AHon8QdAWDoV/yxv3gwLa0krmSFQr8XQJafD2nppA2BrzDlJKpec
C9wqm0EpA64v6akm8PsgvFyxHfGIafQSbTdtvOLSx9bVAMrZCDABmPMU3GBnvblw
qqnlovgIHCNjgfvMc6NkKLy/1kU+hGB+xcO+vdMnKSADSiegVzk/OQRNKiA/hd2o
PbkFEiEO+J2/zeLXx4fBQn5fn+3JsHWowuBdSx4NE8dcRsU3RP1MeE/2rLUZYSOK
bGMduWJoiO0QdxIb+eAPFHla2u1l5HZaYy86Sfyj7QdKxHO51DoB5qRgPbxg/iNT
jhJfSYzA2iw87izfySpfBLZS/oWtB/fLWcIwsk8QSf3Wd9TY9GIHhxYz7RseaX3x
fahCRDqWY0JsK9chuH1J5q0gWl3rlscSOaL04mPHBjnxaBqv1YnKzT4JpANlQMRG
+JXWyvyONyZXs3NirwQ5RJdhOsxyzcBbMhmlC2/xPge5Neg03U48LQh1v7/kygRy
jkXLdGC5uV96Q/u++1c5mOO1SvwZ3RtfLA4770IcMEg/iHAHkcUBmRmZhuGeJ+Up
k1p8LErfDFvElA9scDb1hcapsx1p7P2/xbKTVLOBo5i4G01ySLgXNj9FV5kBwy9J
yXEu51osCDEwIVv9W4+BGgGYr1s5pg8JqqBCfWQkYXBcTG7GTn0S2fwbLlgP7/PW
RimgA+ytYEjBRk9lViMqBaoh+FvpElTKMCB7fZz0r8svE48ApwPJj9opNzty0npN
yczvlVYYA9GFg+eh+IJhlZrlcklVqXchUK3EGf8iwzCCBfL/4EgTZAtz7VlYpGct
xO/mFhTjEaX19Yz0iaenXSdzlkmdF9bZe2GumPffzgndr1hrYvwbHvOiYHNYBNsc
b4bVB2hwG+fsqMWHhqTI+2aAuZz0CuzjF/STqPut7UY9CyaPeuux1Rono0Gl/4ON
wwlo009ViSQBZrtNhiIRExOweEjZ2dJmJKxEIjq4nJgpUycxHmBx7zhBvItHjMco
VPZAYsQFpbtmHPcNLN2JH0Bp5oU3VMb16cVVxYzpX3SnNrUy72bjS5gBgZSxRVj7
Wu9Q6BgqYmvN4YyxNaIL8HZP9YyplXpQEEWh3sOH7bmf8trcz3F+ryU7uG4dDeJf
kr4khc/Qz5DvGzNYGsItaeTSOldoDp/Hy+kKQ12YIJ1eW+BbSQqFD17rVwrA6hAI
XYsRJmTzat+Q5WsmjTbbDMfU72HVBTVQWQ5lGTzn3Pv/PvdG/cbJZReqeaVifiw8
7sDmDBc78kwhXLDncEMeGIugosdqRJM5OwDIP5hAmcvG+lIxX5xdzq0mgxiwhKEg
rwaVRnmffAX7oSvoCaMJEowEW1Dh9Z4+On4CjE4/3O4QKwTOEAEguTrLZqiTdjqK
CD8uX3jlVbanIMxc5iTtePuebZyGl9SWNSRsbJgHIc+DSmC7M9mxT7Kt3lmGjTDG
DV1coHodNgFpEqnCoj2LpwKEZcupBYGpo5OCNITLl9mx8/Nq0u3WsqExjYxixV1y
YLD4cSy+O3qvidxBODt9AeWJX0NVEKHb1XvyC9U7xkzol3R2IGyP9bgukSQueuQi
11Qk2n4QWvQRQebrmrPvRG05uRfwXpFvxHDxhbi0OZZ9E1TWDuvYP68l/iMplnPB
dfScAZmwIu3yMIDtnJOd7BdkV04ZSjFb2h//iXMEAtOUhM1GEAkdpEorjga1MUze
w78yQAFnD8vG+HRJN1VZiFKG84ljw6SjxiUaUcxXmSZczVst1+67V9TL4jBNgdCR
HHeGjWlraV7pmkrZWgS2VzYmrtJUgVULZ7VGnQx3Xmi04hO/E6eexR9oaFMthLOg
4TiyCZ9pMlwkb8M0Nt8z/WUTZqO5ymrl6HLX1Ac2sOTkVKQ4xBtuWnXjJQUwUn8j
blRJ5MzqZB8EPVdo4M8Gp08IU1jDgFOa4yGrnx9fDgvBi5T2tr6Sp6i9ancJv09F
WMAiujJ2wwU97WZYVQ7bAlZV9OIcgeuggqq+heIy6czwRu95lG1TUK0vatKwIlII
01IcZpbyBdoXIxqVOR+xC8IJcIOIdp8QjJhvsRWD4B1riS4YGWKkYGpoWXFKRpVW
41eNBGNKPTA0NTpRvjAWnzV6KFMNfbzshjMo6F5u4WnsHgM5PdPvb6Akdvrgpf/d
PQQ0GlIkpneI5cna0OsP+Pnov0e2jK/jNMKmQpuUjERzO5aXQ6uI9foNyvMLR4GW
fo+BEKwnDBANNMN+09oX2Ykb8LzFC0Bay2wVzfN8cz9fwW9uv2atqbz6V7mk0nOH
rRQLIAkRx4Xm4rivl2pqRnNhKWVcr6TaaB6bC7LWtSmQU0Iir92OdtUoBwheMt6A
uDhklRBAKWeUPy9/hgleL4ttF04t4gI066ppUjXEZH0fSSpQcCYKV/KI+48Kg9aW
LyzfTOHPjQaQB0AF5VtCOAmzLW8R6fcK6UCq2qenK4SU2FzBEEV9owJu9PNcYASE
MVobuX10B8MbYNGsbayzdnxemez1J5NzPSX9tjH6HV5jDttwfqwE7gpSOL7dRC5n
W6YI+KwJsbtVZ6TW+eloPdgWmtKT3ofvC5MWXXwCit9TSS703Tv5KupqmvoOf5mG
4ZKNr62rnv11TkqDA1tEObq+Y7Sz7jBPgCR8HbMdMCbNeJpJmFhQru0EJIkNipry
wN7xWjwQdwas6s70P3cXlDt7DQUDIR++5fWO7EoreWwEJ4vlEHx6BmilPowipC9Y
1UIBW7nwB48c8PvOgj1caQH/EpSKaG3Bb9+OcgNmia6bfdflsUh4Q3+pOPitULNi
LW0ymptAHkee9+vR1qioZdCIkN1I/Rd7J6K8caP1A84GeRGxth8y069a4uFM3lVF
XmyKvsg/A6O/28b8ZknYG8ZuPn9cYeCORDvEQyayx+cZhVGspqStQTdcrMgnuj3N
B7wWRl7NUVnZxJ5RD5viN8jVL0v2Lhm0X/akCgnrSTEh+DNlS8CiMSNU4OJ6u12h
I8AYh7p/xVL0siC1H+UrQZmCL1THiNFI7voHAzQ0B1ROnJw9lt3suT90dvx5gWAC
3Ol3Wyd9JlQyMb0rO0RRehRTBxG9G9AHbx+RlRPaoQAlYf/O+XDilULx01PtslcS
`protect END_PROTECTED
