`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OnzMLwvqqJwpNOfpgdJYeZ0dF4969KeLqfXyOHEZmqrOjr1zfYPkgLmSwB3H3TZm
ksN1ypg9oPnZyoocquZLn//CW0AIojttWXXgdIHjGXO95BqznabE69lNQ4dKZDoB
wUfe91ax69MQlsow9Ez9PcG5UE8YzY5SxetA7QpMcJ+wNMjH0T/9Fqhd3ulUmFXv
YzrDMt6syPcpeMxHvOcM/INRapWBhQEn6ylgJx92BnYZRlqUgJ/dnyqEB0nK6yTD
+GwvJwzOTOoHZwkuNYF4cMEf/1hh/wl9g9N72ESMCTknI+QNfB21Hh43ANTDAWiA
1h8V+r15QCAYmjIwCx5YkDbShzUwEIRdihd8xSlzkIcVh14iM8O2QNInCUJth8AF
hWa/Kg+U4Fg0zxUEXq9XXbxnC7Wzg6HHEidztBG3a17cuV9AZD2cUQUlheEtZRL0
s3hy9d4JWjSVbGWu6edUArIS9gNFGf2j0Ps39Xhdufb1+e1RJGueW3TTQ+L7kNjt
p9Y/+6lrW7Sy7Qj4gR+PTnzsee1hPkbHUJmniAYUaaK2iHDv22Y/Vtcs7qD10eYL
jKl0pcHTYApds/9twQnYIdEj8XWFkLjqEC+bSI2lJueVa+YvUSPo45fbWVhALmw5
peDdfCPqZUZSnBTTQ99I89bZIKtWv6KNcJv9GSaQKO+52+r99MxowKj7Nc4dHiW5
is9gtj0YML8YoCROLTKcg6yeNldSoVjf2dxAS7bM8vDbI8cU2IWEdTYWUb+UodZp
UgXIpg9pBaw7w1dTeaGrOeLtDi2gtKKBfm1yCTOOBaL0xqAU2ibqtCQL3uXBp2a8
Xi0b5bIRskPJvORZoOJSGEqndDpT2ht+RbQeMCUTlHeChtIePfAPapOXDPbDcfbI
CZECo74L/rfBElb/UAi7w42RzRq6VlgtOUe1tvoGug6C6GywppmZUQWNBhu4iopI
yiPiq3b8f0pbjsE2OMqfwVJl+Vyxnc76NuyfF6vS3tpqzkrD2zUm9V5DEEsj36OU
ADIUoEx+Z7brPluB8lhTshRr1NrPFHFrysA49qqOPWsPKhmfiC20dv/UBjyGSHxc
IYmLzjCppjDpp9kRwi/7i823Z8CGDLDH/8W7UyNXL4cYsHtgvYBVVqyDZUKuAxj+
UkVkwoQHAG9XxjurAyIIDd+epXcCv1efEbeQwWatukPtn6RJyBLUEzcZWjE9o7Qx
uKCp8T+JI8ShMjm2nRvUqj6p7tAVN5C6oFJjI8YOlogstIdlts2ncgE4g7wq9iGF
NgLiBlZlDJqGjlXwPd3Z3sXsW587xq9ER5PL0ZuBuDbA+mkSRtgDj4IUtlRcinr0
7TnAe2IJo62wvmuFtxtH8KY9h9G95oShznYVWz34ERwHFPm2gz/r1opFre6PWMGo
uikgdHO6YMiOECTe2ThwEAp10XucHYjonuFzat4XYZwl9GlQp+sgz4MAnqxlfIQE
7y+ZgAlf3giSv8dPn9UuuwRZ8chiYanLQsb2j7trIWBjDyFKHZVGqk3duF4/z8jY
4VqiUk5pK/Hl9UoGdBKD3UwoTJtbvBrcmUXvn2Zy07x0vJBw+an+FQdP4SwBb/Xo
vBQ0rKnw1Qvnnc1pAEb8qWO+oL9YD0CWL/j9Tm2vnRNtYNn3Nyi87thA+K1HRnB8
Ppy8LiPbQasWDIAanRBZ2GwsikqmvUtdbzhzAT+lkY939V/sK5CmH4KcduZnho4Z
yZznIJ7MNKBGJ+WxgW945xDboWUFlJ3KpD1wez2ZDuFeVrwUoDeiaaOdrQlLBY/K
BKDeIL5kIQiF6if84p1v0+fnXI/o41g4b4f1U9mdT25kgzXuMv5mK82VqHRUXk9E
sj3g/t/XTiW2gmie/YZVFNnsQOd8AzN4qyz0ugNd8wyFxTmw94GGWqwjRO3wiGnf
jnh/mYo7i5baaNlKDN04Fs+xcQXXMHmx/GnTKzIC3PD1axv1K0iirgKtDowhgJpx
LCDd/MpcBy+lfNTdoAvhVm5v01eNXQceW6HsS8SwciVNBfqL1ZU8EPrGjW2+TNBM
wNO200RGdoVrK+Cx4iFl2qKQYQupHF4EVtM8o2aNTDK10FUa3Mh9YRhuGkUs8xB6
zHSsBFPhXc6KE1VXwDPOhsA2zZ/tfI5N3QpGWjQVyQdeTb7drt474JttUj1qXytl
kO/ZMUso1M1iM2rh/7gd4JZvMKas3u0OkzYycs8vrqc9x+a25uMbL25X4UinRnQC
aaFhtoFFhJln2D+TeYV3Qdxg1/ByGugj2PxkkRKHy22GSQzUg3FJ6GiBZbILwA2J
Wo65Z2Lk89L6xSMyDgj3S/bVxeLZiLX2m0GyQ1d2BjXtzVXyEJacjdsAabcdrCRv
Y0O4A4AgboF9TfwC55hd+MZW8hUSCxmsZwkwlbudxNZb0N+JIGVuG3eCenuKa4YM
3EpdzG8x35JZBYBcg8NTT5zyxtgGbhPH+cqusUfxCq6rvzOqzFjZJE49le0kSGkr
zHD5jqI5uvx4pUfBqFzr2v84Q/GNDmc9QHzkB0C93HRGc1RjWr+TRpnZVDMMoVj4
NLQ1nuAbf5F/7gVX+hdA52DQ+cRpwAqjcacP/khRW+KAiludk3Qac1nnvXbDNyjH
8/8as6byXxRLLVfODYL0qn7R5Uxn4Oh2mbIdN7tRXhgO0u/fz5OVU+smlvAQ3BJg
OtP3sNU2mBs+DqEhqFNGwtpT4fdVhwG/bFlfhySAz/5J+2Fs6N5jK17wRkNmo5AO
Y9EKbS5Q9mHJpNo2ndBV6UjCB7XOpip46DNo/wP3ro98CoxBj5YK2/UT579CdKSP
xZEOqf6j5Fyr9PaKJ2FhvZB6md5maCco8Nu4waZX4WpSqCRntF1QyGiy5xyKiiRO
/kHcpKvgjfq8deJ2y3ubmg==
`protect END_PROTECTED
