`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkzbTIIJfUPhfft7bFXyeVKIUv76I7cYQKQq0Xzl89E3+if9dv8YAJrPUe9f/4sq
RLR1K/2bMDlYVdJstWhOZa4qU3D13dy240ifkV3WIMZMEfoZ/9v5fb2ILlA/yGDp
rA/SBJAwXvUuTUa+PtMBKiI7nkFqg29G2URTP5fes7FAvU3Nvf52qH2Zk2YjY85O
j0hV2h/mQR+xtQJuJwXzKwGa5OXW8pWIO4mFfVjYZ/bZWw2+RN5pifURKpfw8c5+
gT3xJRtaaMfsuc5NxqAKyeNqoIwRqnzG1uMwWrqTj2RVOjdhvTpkQpUIwgGqIeke
OuBDcnlQr4s/XaYFQYY83zxSSBak++MeD+CCBf8QkBLNbDiR1XcTig9h3B3Y9Qxa
RJKsmkt9jRIu8+Fa66lJ4F3VANnXnBpgglnm441Q/XohEcvoJkyuRUiBqR+BN+X0
4k8ySZ8zoWLbNYvqEqDGnw5a2vFmoGWZvaIhSuEaK8EG8WXQGQSmlPUR07PIXcp7
abMNxxFpKGyyrxfnV8mc+M4ShKiLWL7BzTdzekTuoU+rV66QWPI024GrE8K1w8nt
8Ozc/OTnpq0lPp1kk22dPIu/bfb+Ynd08PdRCE7s9BUTyDwRsDl/7cw/VhpUXH+T
zd/c4q4R+bvhBY+/Y22MZ6oAkyDZkK1gCnboU65w3stAUQRigyKr+1HSpYejzf5w
ys/nXb0fp8LJJQVcNoREAQoUiPq89Lawu2x909wSkzBiZbsNqUUYmXCDfr9YlE8v
52c4h/BSEr/7GCjJPOpq2U9Op8grszF34zMfb7v53NCqPJa8mTqB6uBdoDtbpTGu
eKKO0xmS1Wf9RJv7amVw8z4mmzFy2UxXmKNWUXnfUyW0T9Szs14DJFGdmVI4tlCd
evwGexVBZTofRAmAVAiQJKkBqHwhmBr/cKh8rynEgwgYNXLTAkn9tn73i/sg7pYO
E/qe5i6M5jMYUjlrotXvOyBV0EDnsVKaVwhMyy92ua9oSgLNokzAQYPALB61TsoD
+pMx88DcIQtNqt4zNr46DVuaJKGfTbaBCv570FTZyiyKzSVrTelmE1iZMlasFdPw
v680RUCwVc11LKjMvlYJbnXNc0w6fuJfvvjrju7OW1HQ3KTxitI6baq4fmDqn3bR
u++Ttw4Tpn9daUNiQJLSTi+BtFyxsE+5cIup5/RXZsTKicO6BqsD7qsqmjlq/l/2
Ttaw31Y2Z0SWlG3LMsoNuJ4pazgsXc6au8KCeueOAy7aUu5AwIbX3ENKs2kiZvJf
6scp4xG6sqpjgRkCr5OgN9eWNLQNGLBLCLktZ3UicFMSAXwlHh3iK53cMJpw9Cg/
OTOgcCq8dVaXvcSO+F3eRLbbEDj3n7WR0NGlErgXLxUzRv3fdfnXR5FLzRSoGoNM
pbGRhDUASnBUEsNxWGiVugliN+FSi2B/18n7C51yTB36iM4MP1/81CEqxFuYhN+H
TxVgycB52joYbACIYRs10HesQyWvFkUgFl4I9Q2a7bPLSBGglKWuQ8dQSE20sHMl
CYIvrTD1EqR4lLiPFBWJdXaLVDbdAWyLVxqEyimoDcz4JPMKMtqbk58RP1Vx9rw3
HqhKmL4HyzWhRITL+uFb0rTkRtQ28LBVsz4/R8SepnMOCB/MbBr8tdG30fUBdNgn
GwYS5l7hjhyZ0TuN3UNcD/aM8Fn4ZsrIKNXC8kHl8gSFkH76NvCWAtDX3vZBQ2oC
LeHKmuQpDBm0FySCtz8cgyubk7H7elzNVjho4NeDTj6ri7lBbXf0HtmKFm1RfjPr
UOqjxVhZaalV/l8n6yACH3BSnPaTW/bkovcCmxXBHhi4kDbslp+RAksAREslIYk+
5Rh0hjRmp9VzaW5LSuIBNjwftWWIVqHF0XlX0vWc9//5TItPVHkonSO6S5NlNXmk
Yai96Q9SEROe81gbvc0bYDqdaF5cfwZSSkTr8GH7D7LiilbEc4+48i9D6+nPmE9z
UK7BGGb3wiqYrj0afSPZPiVcUVk6xtV8/Stl3vZP3xiEXyZyWwxT/DXcOYS53bm3
pIhclC5lF6bST++OrKTFLIs0LSC+oubBt7xzuDQk7s6M3WXkJNA+Wa+NMT7apD3g
z+Vk5LCH7E2+Efsr2qt+8mH4ORfNmMWnj1j0XX1drcL0icOQJ9en507njL1/kLlq
qLpVD7SKcI/l+dqLtAmHGKZGCWHcQJDEQK9lUbQkYTk3mGkxmJA6g4XRL5vrTyBh
5LCIvOGVFUb1LCDxuSVxKy596lpkMgcDnKDqYjZ6XX+QRYKtVZ1Z7x4lz0B/zosx
Ew+MlfZcdj+5YcipHQ3cshH8s8POffF2+bQTBfC8EuR7aoSRW007M4sS5tWScwXB
rn6MxvLwQpAgenP2cHdz2NJETQ+UNvT190SUPQzk3LDLxmXZIJG+Php2E9EqJ9kn
P0msxKMsn1IcF9lYJ3BYuyVG2mOnCwa0TgEF4AYpT2c7clbYZzT2aliSd+4wBhA2
SmPQPX66SfMlb05WI5oDbqG8APjHMqNt9B0qqVGZ3YaCAjyjG8ErRqDfVEnt7WFd
adyCh/43VHzKYlqCkBBXZTXCV0/e+vhxPtGIwmuyakDYQhBI9FMZHW/UYpVME/Wy
CbnbLIkw1KGy8OEZvt1emqissq9zxYcYJIyQp9sGZM2Oei9r2MavANInbGmz0BFn
IcTMVKYe6qwXtSRcm6CmJd60h7VickNCs3RbaAdGf2cRQO8Elv3ULf5/ICXl4MZU
1r9pTs3MkDU11gkrF6KpqAOAIwbq73nRNHRgF+C1pJpMbNsVCq8l0MSrlZS4Po59
RsbNVEmnABmd0Jr9y+BvnKATQomHkEAgmzgCj2da9qkB+DAuMpF/UqMYm5IhRbn2
R/vmyxD11qFhIt6lVE26RiajDM/9aOcJuCArXoSz/aupxLSAAtwyTpfoX/QgWFr9
eELbxo/qfGncRSE/cjKaj+r/KUH8Wvih2aS8kT8KAnQIFg++DPcNMuUDviSxF8H9
craTjlYUuoO0SLzNmv0K7T8djq75GDGu9LdS9g27q62oa/TYHzI2cPjLXNc9sXVV
cTAGTrPwPb8UkCVGnZTZum0BkcUoEgi6rwFtnjsTFuLQ+4tTgcjca85dvS7Vsslm
N0z6a+Rn6fVShHF2D2F8a5A0U+5ii9tzKdmUyzT+bkUoaAQX93L7iyuX/+lpIoBr
Im1G20pP0rZrjASOJ3ztLSwIwORi4NV3pt7ACzb9eHEZYcUk7FfylHjFJJmyhpWv
ZBsI7X/qWFvIyuSNP/ZiOhGVXWVwWIsA/HUm0cWWXi+yL46hA4OC6bSvadhLS+kB
PQbckxrXuAEClM+J41pcRQpGHyTOE7Us946Sdxdm4Pwk8WbO7KNH+jkeNPZc6Hkn
tbgkBxbspHlLrKHLcCq+ULq2xi7afp7QorjnqNGPrakB9FiwASfasc4omzWgHnGM
PzTQKE71WmUPYxvQBcj4R/dnxGWREQBnzcpGh75F6JX+1pdm0tyjUBsXA17KjnZs
uxnaw/8nwmwlBKs0Edt+tjrSj7jvB2jvnFpLUmcFUhZcgO5uFJs8wltDo/fFVWyb
VW7nOykkcB0ZJt3CD9cwIUdrdj6tODx5K/sWuCiss91pJ0FqGVS9YLnCR3A1Qr9e
UednCGVTdh3IOWqwO/k5LnskFLrZNq7NJKvA2f+YwIGhH0VlzApmuv5SRsvQa9Va
U0pf9ZVk9v26DeYQDn1kgYbDvlz4Dfse8U15P3cEPbwmzZKIzpwFRFa6mtB53NjU
Pk2SkOsAfns+ZTMvzI9RVKh37+gIm7Tteuif+B2EAxGtLKlzKrKukkW5fWLCuJPB
TDM6wIX9g68/hyv0Kk7asQ985Ju7CYoacBWhkwcEyvlY6n/rIAGnlKoJwSdU7ZfF
rBEGnpC+LiUZu7w9S+R8WMVQm4oUYQggD5fb7XZe775E5GmpM0A4/fvRBsViWTIZ
M/kpANqFtpB0W/JZDk+8pdC7fboi4t3yaQkJWjSZCNhSeVGLKkd82a5b/bmCn7H3
zW/0CacZ9d1biqiLujNZCPjYM7vCDZZiIOwSUgFqjC14guwdCWlQ7iSoxE2+9mBS
yT6HF6TzBJpADNU1GlEjF461w8FZtVFf1NcjAE9VQLr/u1PoC0YL+6i09pTLWp86
tOh/0PkVF7uEv4d6oTuNUP1T5vcp6RQUmuy1OeuPQKIzmVORkXNCdldxXMDS6mEN
5v3xmUz22Jp5o1Le+eQdG8NjAiLcBqaIOjwun3sSu2Dc/xCy6LYBjZlCnixmWWdB
ashbAYp9KqbrufBcnF6reqZ22mcyWbJk6M1PuT5u9IA+WBgxCXxv7GjtpxAM8V0+
sDgZTbGm0u4gsWREJfQFQNWj6BPR0LU2Z37M6+PwOdveH+bRnOb1SO2rs+t1JpJa
qBvObo+IKv5z7Xzi2LDJ9fdJwm4XSnqP8HTci+yMHaOYiUkxIIjPzy3AOWtPjf2L
OpGR7dnqgQ0/hH30C1tWnCivuX8jvJK5GHiN4BowjJqcbQs4Uz01yC+hEfJeLIOd
f+x4K700WX02m1EJEWTakySU5Fg4eP4kriuwK/exOEnFXe1s2QfV6/It0ZmL24fK
DZLCZh4rn8KJcGnXWf+2nLBcqitHBe5hw19rLi5V36R5ii8Sx5kgFhR7KItAdOoE
IrCNZ9ozUhUPKkziZbH3Txx+Wack1ml9sSakImt3qjJSmP69si1LerN2BEAgo0Ln
uMCV0GjmQI6BkUPnJQ/Kbb9f3HILxj+ET2zU/4ia4AhmzRki7h27tRpPU7u8HIeq
anufEM5V2O2EI6h36usIakQHpPMvl5VHyMgf+haq6hsNbqUeLUs9T9d+UtVn1yrt
RG6FgDs6qXZBTdl3CAFVAsgRwUYjnG4XmLXiMX/R+EbYCeJ2Ae/PrddBFi8eeQOJ
Ojn6tQDDnld4oPBXOBC8uTrpKjNkpRL+Ubnca69X/OcJx4jRf38WjV6Ul3Nz68tc
Ij+PimbxjyRSeky2Gew45hHXPANHyW12+vd4DFPAM/3b9vjEJ1ZGll9WzUZB/rhm
ElVXWimv9aEFHWQGNJUmvq+yuIVwCl0pZP/KR1sH9OaKfKLAUm5x6UT10GvaRl/0
MqR1WAE3Ifp58Oakb/5wkcCMpoXunX3Cv1L3+mXluEL0typGex0zc7TMdSdAWayX
GqBMGDINvYeFi0zBxvs6pSRwUOqKT5s+kdagGCIbuDWN6QlcRwADq5S3SfJzcm0O
SHraxS7lLqndhMBwxYR1zj28HIvoEem+wGwDS3sSRqHtgXzXEH1ujwYYCRjNnnTu
ozRxdJfysqlWHIoJCdEJFbdqoD1/ndAS4p/2FnlZNmSt631veqDb3Ftt7rnip4DK
Qr+PDiYdcmZ1wVrfTsGAGZlsTLM4FhthY4nGd0aKbzyDFkFOeEeeAMA3hP67aFLJ
GSnIFVIxm1sPXMQlF0iC09OZDLI94HW0gepwr5+Meo4=
`protect END_PROTECTED
