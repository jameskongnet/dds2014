`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gR2LSgWj616e94QwfMMSzHeKftuGsF0C8oktLLdrdVoF7z10I3trMq0G+RkFF2UN
xT7x2XxOkBgGL5YO/qo0CDUsZUD0HzZTyz6tOsSQKRp7noY9dGLE9LduHCkhS6J2
brosRwhp18GTCpzmRVDREqfr4rtEt/9tPEXh7BGJhMagosrcHaMR4nB8fiI7rLrS
aoMykBZB0tZQYA1uUHBf7Qd7WzgOmNs0vXvlDcCp5J9DuckmC7HBhGYq0EZDqSDW
RnmawyUMGoIzlT+QdT9rOg41BPeNAzlEzg90gmGQ+xM3uPvNKmF57VMuAAXQLVfo
OBXW/ECSlwWdkijQrHbJj0wQe5+Vm0mt9rEYJSsjrWL/Bksywplia9MOKyc8O21q
KR6wDN51o0oqrL+hSIHALQJlFPubc+dW+aqEgstGamHNM1hRU7JGC6qB0tmX3NB0
TbX0JaZlxu2QkvneN6reZptM7JzM+jl5QrGY61QJJg44OpSZ6AXUg77fBxPH+lG/
8SrCbVRZ6CpJXH3evK0/ncM4wiwjtsdJLtE+j8grBHLunDP5+I3siD/GQkojF6sV
/1RkjmIR8o9EVHHG6kwbf73EAsdz9NVxri6D1kC2iYfsY1sNeRlxp28CBQ5UBzF7
SFw+tWaTdZ/XTPqAApxRPoY6O92FMxjQKqLg80nPR2LfcT9AB+CTu9uTxUFamwnl
hMbNsipxndIOheMjtt6JVRHfoVu8ytmgjEwDsqbkvOkdMRYYWt16gZ+G6uj1p/tK
u21jcJVbfooS9e5ly0DqgZb9C4Qrm7gnxcnWJevxAqKlifHs4BkboiE33jaebCmn
F8c44/WxYeHZwgR59XsgdcLNPHNgvJfoPHxXKD/igYmrAQpAO0Tbl3ExyG0vAsTg
SAwEk5mWVGpH9frB1Tg6o79VQuAgLH9YOePCeLBSR31jF2Db49v19YDSyL5yHbaH
Tyehsz2d3Vbdr1hStsde3KzLqsLqEkGXlAiA4ge0swkqtTpvl9LtG6tKLHxAnh38
NE3uAW0BvBuUlUV8GB3JZe9Cnq2WO/en6w66dCRu3GIRfLInLVz0DeKu3huK9aH5
NyBtgEjEB3tQQBoK/DrdB1VucFHOi4nyoteCvGXtKB3NiMt7G4izk3mJmVw8m070
NXyrW+f6av8ozGGUUm3x2TWYES0IQn9IaXOGTHt8kWRIpI09ZYKakpHMZiBXcvju
vFaHPhDGArrKqIkMzzvNDK4RUmZzR64iAdCt67Ba0cBWzZb04da79HoRysxNVMVW
jIAO+HUnNLl5JVKIBdkXQfQk8wN54vm8F0M1y6bblBn1oH0Q4/PErrZ/lUAGqpf1
KJTga7UtALNVzpfdL2GpN52PZ/u87/+XS6e3Wszu3lju0eQWPmTCB1Ai1xNFBLj4
XWfF77uFplNkRLs17IwX5aT5gipjsMRiv/q1YogFUmKNShSgrzJHWck3KgiAaZsk
HBfV+eAgPK1Uc1UCI9VV0uT4zfOadFw5jEsBAxnFXc6mHnAJNT+TbnAEIVPhp1t+
YUU6kOns6+6dcI60gX+DAo9y4U9NZHCKXBzrncn3MJXvf6GhylphnuvrcY5dG6dn
DNhJzsEyJapG3lzJ1J4WByofyoBBOqpSBcP5xlLTwEq7j7RqSBx86WIvQK9gep6k
UUSQoZ+/ACrvFScCFs2LIHNJ8fLf+JMIb8DUjjfBMub5bkIZMlqZWVIFi3NB/n9/
1FBtot2eh6WRoPSCBbF4/fYm3soh/LbiqLMOfyZz7LpJpRfTHo6RNbydGaDe382D
F2UXIcSC0XOaD4+4IQuIVcNJKAmHcptgZlNO9gcmCCqrGtZRopB/NgcQOcjXfznB
nHL22JP+NJeXGyoNHf8ieO8us/TIC87Y0t0MLpgmgCPhcMAqYdSE6TW78PiUXlYV
ycUdqLX+w1H9uL2fc1Zx8fSFmnI1yWh/dOjHZOIIHXl31M8iS0WK7fn13em+Qorw
p5YnZ2UtwdDLYG01hP3YNkoW6kb4bVn46hi3PAHTsritGZ5NitYmhdpBJH3tzTUd
KGLm3aY3DGQZkcwmuQLidh9prlXT54gGZ4Ux0T7stja+9Kg2Ak1IYVa8SYRdY+Kk
KYgb6jk1mep7FlA1cCkWb7WPVLT02Re/Pht4cpjtTI9BOo6CO0q/TNtrNzx4Zkby
DFLZIFMCdUgOL8haXQsAY6p4RCvkkCE1m67n2HPhnz67O4ngsmg3kC9fTbTmKFmU
eOQaKtp5XmbGk3VuOD5NcWltW6rW5jjRaKChwdcZ3EO2J8AZShIl4SIng3Mj+HYO
4x00380HpDCScVqdzy2k94dFCWCGh09pWHRe9CoXIIL+H1Khc8biBQPI6W9MEUTw
TCxRY8s9MRY/+ZXlL7yry+K1UQFbO45VYouIWUCCNN97uQF6dbm2uRxLNlXoyFfN
AbeC9UWw/jMfUTXFrif2PDy8AhwzZ0+FULYl4QZ92Pl3IIHGyXkZypXMCldJxazf
5hRsiWEgk4ahE2bMHEkyjPs6DtpHIs0r5+u11Ft/hOgjTGVn93eVskViixXYUBlW
9oa+dj1vNsFAaADSbZ4tscYseYj9+9QJ9Vubv3SsUYM+P/LwxRUqL6Gga/22TjaH
Ez5akQ/bfxkN8GOrdTC/acPHRD/Dpyf02LkWRmwhxtdNtrDPOGbqNLrwOhRytM4X
rzv7Idmb5cgOcrAD5gNZlfxCcpuHjB32a76yUhWKFzO6fnEdVEZ4tgwgMqkam9mf
QqiENCi79eCNNxv1boNRcEU4xXbrroetiGD0h9Xpap8huLS+h/EnDZsGEg9xx4Cs
IgF40T1Lxxu/rg6Wug4BNCe1fKGzVzpUtmCF4XqfqFSzwOa2Lz2y9645ZrEXh1d2
aIG+FyEGd+2ZujUzIQ7L6oFKbDjpGlAP4V2WA5zw6RznmpfO5A1BRGARnrcF0SMn
OkaR+LXWnXS9f6Vh5XgILc4HjpwwrIpJ+rIY3tXei+UijPKzMxojGO2Z0X6/s+Go
mJ6JdHqfbhcrrBiLIB75dd1j/bQgJLZq8pHTZetva5nO2ucGlLL6G88CqOpH8FLJ
wmuPyYq0HBBXuLCelIhHOFPnkw7DzJwFoK0eEdGDEBjjRGY30eOciDtnwSetZLht
o1Qmj+3D4UuuUBGLjONEHiIKoeGy+LB6Wzeg8rUHIlZgaJSfncxsu5M5UL6F/MnC
Ge7ttZsL0MkZdbj4Jw2iSc2xofx1jnQvRemIZYf54CzG/CYP8NmU60Hw5VyPc+j9
UGLMFmXf0bt9Gyo1MCIERhnQ6VLvQSkKM9HoBUoc4f0gYXuck701XS8vVTgf6SFC
kyezVyRR9us+P5b7+AG7Nn6DxwHVHICN7ye+3LG5rJPc7Zx8UMJvoad6/13TZ2Ih
bp/VJulRQcnUAJW7HVdgP/3wwHKOHmRQXGsZQWj9WHvr2iaX53xeOeRGJzOdjN4H
hwcN4RYuKgu1WloiwSpOAy61qPIxyrSSHCkB5OlcfeXXrByAXDXb/+LOietm/3Qj
ybuAOyJK+/AxtkUs9VfRvfcktwnR1FrrU4YkXB2TmXQ9XNnAGpFLvc3Mgk4B7YDr
jT1Wctsha4xOnygMIb+SFhVdKERUK8VQtTIJUlvactSMPgbxNMRQUqtnk23OLb2+
gZpW2K281bZw5Hw9RxHbYYrZGQrs0sPXCW6+5dFZGwBJxNfSEbfrYmGsCzo5Imxb
g0gjdYwVInANw8nlhA1fOHfIqiwft+c+J3LybaqS/HYehC1MG/rVO8o+e1kMN3hr
ViGxEcfNP99VCMd+UyK/3x4Ur6bE2e/pYhlD0nyhTW3d5EGBaSmUd7x2Epxe4qHq
BSYz8oWgpb2EoKdQOZiqK6Sd2B5ANlOQSU6ibHSDwyX6SSpEN/uLAmsunvrN9aQR
jE2jLANJjrZ8zdAVaYfX7KD8UC7yO7o9sdnX3GvbpKm2ZNLJvejheIa1zNb+cSTP
E3muYxdWdVFiyzhie6dGSk0/5r7D5mxMm8sfFHivmJI=
`protect END_PROTECTED
