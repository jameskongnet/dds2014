`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gy8dEAZkhtjq1qrdo2sQFgJwBp8+cCXS4cq+VWiPCLI462yoFlfo8fMv9kN1/Gj9
ggXgaibHe3LPA5TI6k4+gJC/X90ViIPFsVKDUnQqjRCZhtqlv4YAH9VxwhQRh5Bq
tPuEoOpNhRep5y+I9wzunEgshSxpO1W8a48bTCWmnrB3tYqW95oPe7BogMvFRqzo
aXCsFt7IC2yIwz0sLtfc2TlFznbCb6tr6Nmfy6uuahFJ3P7GAGth9ffJ5w+1biaW
r03NNcAbkzfOCKezQQ4HW/hPTdia70I2fG93ktRMWWSXXCU38j1H/OqLM3Vzvn7T
KUG4v17H0LhyA9mZmvH9KCsk2kBpYLlzqHYgzkeXB/V0/4I0IytXM92p8ZMX5H5v
7As0RnNSRm8SO5eG+pQ65Pfre+hUafYScH19dI65pLeoLlzsH/A5oeUf9gY6KZdP
M+tMkJqLBONMYDSd8TUJY9KBnizPJCjEuiIbOfcUX0tkYz5kTQ/5DdCFk+vFvREz
yks4JVV2sPZpLul3zTeeVyph3+TI0mvELEffHy9Gj/CDUCBSoSwBhTrU/cHIo90c
YJKOXUimqonmd8Q9/ozorpmyPVCkHa/+aXzdgwbWuQ+uvOsCm4CUzoIqdJWLQw47
i2ozwWQkl9D87dKFCBJNavVVcaJQ76l1NLj2BLiQ4vxSwskL29+57a+os3NZf7qt
MsjmrZfwVbc9x0tLyQbIjcxR2IBgA2ZasdKeG+BeyxwZM4kx8AaLFHuk6Qt6n3Ef
a6UWJ2gI9QxLxfN2lcbf9RkgPVaVDg1rwXd+8gM4OiaoQfpM4lbSnPR8bJi1sUb4
8kvVlR51I1yB6y2SlG80k8QSM/qonVysVTTEWJ+eSB8nTXJFSWcrPNeO0nelYY6X
z/649y0yAXTxHo1swBPzIaoX/3H2jWYrqT0Q1QBqzSAnGNaHpfQJFepVq+JJIIGk
54oirhPW6YdYMeECZ4QrHuj5nOIH4Pkzf86zJgPe02OM7qMLdPPK2vXX+KsLFhLo
9utv/9h32JC8zx8ZF0spSpCiCnxZhlRUSp4+pHe9L+TvFbrgqhIWSkGs+EfQFEqr
kYpU2GuJlgC5y/2yE5/XfHkXT1XxCkhiSwBjz9IX0satV/3NYtXEzGhihNLBVhe+
6k9hfzimJNzJZ2Ge+9ueWn9ZLk1lwZmB9Y9QefLPETTBZ5yuzjRcS6jxiJgRcjJL
JqBuxAaVxFhGhEranxqTHnd9ALUYiwOisEFi+5wHmsdxS4tYJkxeiOOXads/12kR
rzroYMI9OAIXvK7U4Y/EJFeKr4+8TsksCs2l+d3Y1gHCCANJWhu7fxANpUflrYGe
FhioSD/a+7NYORls8ihWvTzvj8FLcmwZgut9l3DkVENXFWZXcskLXEFdqGz03T8a
ZA4RfAAkD3kxKJsAciUg7tmdalAK5oe4lovjkWAnjz2SiJ5rymCbW4HRh/3/UjuX
oEYR59LMMD9V2LlDchDK0GtDjQtPieFHQihuWm4dcdk=
`protect END_PROTECTED
