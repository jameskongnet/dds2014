`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5qcJLybUBrBsDqYOeu5JVb48LuRMSV1wSvAYH7HrqcC+jT2w6vUZjnzp2Rc9y83S
4pT/bZ65VzXQ1/cnQO6JxS0uM5YNFnwpJGMiJCpaH2gPeRSNwX+vQO/RhIluFmxg
niOT8idnz20MGU0oKsSzlh2VFAqMr0LuPCmq9j81Wul/+gAYw6Q2RKomizb5ZKMV
Je0rTiNi+l3LrIaIktgbmmrk7oScjQNwmzR7Ynp8eTxYZqM9ua536fk1D/KQvwfN
r2RaUYpkV4GpZ2ICqTZkAj/N+nKgFp1I+fF61WRunX9RIvypKDew4xHnirvdZUo3
2AAz71JMte7UPglHeAtxWDtqusXSNCr5BiqQDrfdCsL8zxa9tcrQ898CboGM8hus
Oubxwfsuhs/Nr6nagGuHaqecQmLPBz+3DwyKFsPvy87ABnZPhwZJWMOLsLWr8xrU
WFtsB3doAmPETfefVv4Hd8dFhPPDHfI3IdtjexrT3fRB9h1puQ5Oya80XsO0ZM1u
PmDwTuxfUZaxZ5sn3jVtWYRzLR1o0lQPfESiMzmnEA3hoiE1Aw6khWECm6CR2lQi
XTk4c8rfdE3Q4Z8vJfzKRJN7A5NG/k7ZKDu0E2S8Q78cagurh0nUa6jnnrgo6fHf
X7WZkm/4jtrZ6QOJrp/yO/X4jhGzA6ccTKBSxiizGhrLMAl5XDjCZ6FVDs11siUB
P7lWz69CeJulh/hs5k0/AzaXodwYWFGpBfyPHpZEtSDkNURpJYn+jpj4keTX1kWd
F219s5hfxP/D0jY0y2KPpywmN2lBPpGZSPJfwJVtkwkFHOwxaNmHf08daoKHr6Di
cPZDq4CD0bQBqDdVO74tpP4EQeCBqFXufhNPnaaEOEOoTLzeOG5NuFWwrcmlwjkm
JSHd9TSS1/21wxWWuksZnO3rHf3hEqlPvWm3EEJMsz0n5X51W9yocX71hbJoS2Ii
SWuSEA66helKYElu0oU8BPdsjbcRsHnRX/hw36Ydoeou0muzrygdeYK4EYIzNmC3
BDycL3MbOTOSRAxxIrDG3of+qQfsfp8xj2VEs1qO1ygoZ0pFpZWio9TKiTVan55L
LLwLvD/RVF1P1yz6gkEhnDmvddlRJz03rkV7+6Mqk4OdAaezVN/7/pANOuRQl1k9
AwToXcgjwvzc/Wxu1zstZIrRuOMcnCxF6s18T0kG6A8qH/19ABjwRWhZB1Pn8ChH
jFpMFTgLuiCVZwB4lrgCOt4nK+iJ5jWcVvSHgUBm5XbyKd7/WNqbZfHDZCkO4VEx
PQB5sw8szLpqo91jtpwaW6gi6R6lCJJrGLqVY/m5lA1N5qNGPge+9hMDjYAwRFZt
B1AMxVFhedKa8PIkyujDDptpxlcIGXfeR/sxT09wqG1SyGBj746A+GDAJ+v/3EF1
RCbbPow7P5EN9q6n56w3iW9rzsFPJafJXh0OtJ4rr7tFfI7Y5Amxlg4oWKiFdAN5
onqbPQlSVE5ebE8IhLT6FypT6sXG2J3Q9AECPCgSqMfTv0jiJLBqa62/2U77DJAq
zHMVh5/VbeNk/t3QDWtZALCTdakYBTvkz+lzEhv3YkhJg+Sh9HGnAkLOn5jvbxiU
BWqkylPqYBmz4NMCQBbiKmw7OvNjwvVkdJzxrWvHEXbjoJrCJ0M+HXjJoMn77toC
8Y/WgsRSOlUFTzxp9r110T2nBMu1jS8ZqKs4Ws0DFYwP3BevKkmabYjgioanBolZ
ss8p+MElwXPv60syZ0SHj3Y7RPusR/pD+EM/hQM1OMADMbcdYOnWyqIswFrcUos+
EDxfrfyOE12ENSeX40+1GViORt0Vytki9ipxu+yg/y5z4eAPstoF0ASQLkQJcYHs
uvYZuc5hUjueIvOEE+0q+ja7J47EL03V+W6ujvfQrvLC+T1vFTE9FJ8GFJPGBxnt
SlSg6dXrwYK1wA10o/WOQNiPvkZDnvORto8VoCuthGIQdECuSrDRCXpGLm7tngNr
pKOElOBba5AlTe5lKZhxsWwnPJxep0roi+HjVCIvqsiPWrcDl+8VxRh1B5q8K5Vm
gFfhP4hAIcExoGyqRmtkjG+IjYe75V2kWY0BXO2KlPhuGh4/tJ5Ghw4+3z9ZHXeu
PYv0nvpYWq66sTNchNXUw2iEgKFn2fS58Z8GoeZHXEiD3pVNs78C/33tPVb6p7yn
d+Bv/T1JknFDMV1yE7dibELDV4kzl8ZCFYU6+v7OYAFEX8LtQn9vWvcFmJ12rzgD
T45pVjOng+xTW5IpTO0TlMiDw+dkhB89qJfZ9d3q7MHefpMT6bWiNAbgzIGLmQ47
eF5EtIhW/klFQzOSoqFm+Qx/ZAssJsSL9yKyMYNvI0Hc06j/nlJUzvV9a4MSKxG+
dgb0iDtc9JQO7XdsUTVd6Evt3eTTZNd+3Y0OblAbqEOJxEwRqXfnmFvxLceus6yC
s8F5bvOhVryHTsX5VxeLGny6jNftYYlN8VHOKikfn1ddDLRyXXLGkgGXuSN0spu2
oJzSN3C60M9mNNZ1gVMZac4HzOydNGSZwssrFGyAJwfSt23ewmb/rCcaGm9Dd8ZH
o1s8NjQxQm9nIEY5MYZAfjpp0PAtnD8En9WwdGodnnY+ImcGwzmdtrvC6fnlTgil
qG7A349Qxo399YbNoOrAlfjFplTU86SX8DtPYfSNXZlXGDfQ/8MHb/tLFBVGRckw
yp03RoEuuNv8u/UwEcb/aoECM5gG7mK3Z71+/7dKgmJU+/qbSzb9BCRBbgdIvg+3
0IceeLtg3BsL7GcjB98U3Rjqmk+bFCKkl4le40Y9qv9WZdIAfPWl5xjktTBIEttF
W3RgnikJYhCt46gE0DKtlBeBN0WpSwNvUIDBAxMjXuGbJftF06Zr1PCSVEBvkgLn
Wx70LCLZTTP50yKMJ+E+bN1DsLPzCEJYXqQiGKn64RWBfnAA5086mZVzo7LdiHh6
90KszgbXVc8/ujRyHSa+JFhn+JIv6zftHen2bsaQDaUMtXCbNJqi5CKS/EfR436E
psSDxOYytgmS++eWzEIp5BKSUD+BgZPJP0y+mg6BP/SypVb372s0Aa2hKSbxERgh
6MPm2YNGb1hShj6qAcWRnnS126LJjAIYgdJ3wcCNjHtPQWds+UhciK+eptUDTBRK
y7Y4j9YPPMSAKy9RIrX4AzF7tLivjq6wsWVnOkHH6x+OakOv2Sl3SMnNmsvQUELd
RycAEYxGkbLIyZQgQfQyhSEeXLb0aJ4sDhE8QjtgNG8vlO3ntSpoMqdNJ74HdUK5
tjORcunInxwezOqxLub4r9of15UUgJeO20rClFgb804kNXNedvuT72BqeoH13GB2
pbfk5WFkPySflwyfXxhyUQDuN/xJByORgW98AbjLEySAWHSyMHkE0d9wVexWn9e2
MP+UaVRi+05yqG05V8NFMCwgFvkib26hnvJTdn0+6SQ=
`protect END_PROTECTED
