`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qg98ookmgsY+YBriG6S2AQL9e8c38frDYWAk+UibcjYYxRRiVmq5v8lEMSo1Mo0Z
/uanwD9EackQd/hIfz7VquyWq6ePMs8/gAh49oDBcHssFVYNiqG1pV7KXLKu/QB2
dShAJpyGP8P9GLJ2igsH3biDVPUan5FFdp0cGa8Sjv1MJt8R/NWpgLGBG2WTTp+s
81X6Q0ZIvEw+SB1IBL9HcqCw1rLHNYnFG8axC2bLt3ezne3s8ajBcOHe7wn8DKfv
06g3YNJiFWTM8o7YD9TNWX37Ecqcldh9n0+hjzvk7x/cHPt4E6IkQami/a3Bqxe8
ELDcPPDZRkFUO1sMJOoG6q6yXJVhpV7M2nRXkzyVeyyxoJtQPx4hVB91nFMTrKYJ
16wdQCvLRQ8XXGyqlNb5M/ywt9/dHmISAHsyxvk1iZUBiBKVdWIKZdTHUv1QF2rv
u+XNb11K0vUQbiAtGSsmX2WAVY+e9gDG2yMLixdFYS7Dvz8Yj3Sqh6LR4GlqApxN
cfwpLsh3A2cMR9Hq4vfTFMHENRCt8p6XV2fymXjMLvyKxxB0GLSTzdStAxe4rYiV
790busWILhovQSqsByA7itdQnbeZddIyE12ZH+AqMDS3vIduGzmvQdOPLkZb5bfj
6T9rXt3h19UcV8lS7pcgNn4icOHkLKWzh0kxejbz0GRhCXTz5pbtEyTutosjTHm/
Der0dD9Z14/9iS6+dtoYWV21yNyaoG5QwpGKEmCmrNo+6u040KMpEPA0xNldxowV
BRcxk+8EQdzlXy3BC+Q/qCLNPTm/gNBcabUicXGJY5mJbEwwgXFe/ML/a/olQwPd
lAhLLerw5X0zaOssxQp43aVnRkKTJinnLcQyJ1wZOBYkjuEOYELuw1xll7kmP20/
s/EMXqOhZB40DAIPaZhetGLluE5xK4+0LqvuvA5dln7tQbI2coVojbUyK2MDhiaF
S5IIjPuldoBl9ZGAh8eyF20C1XaB80/R1h2nTr8CVw0qU/rV5G2s1zpPVwFBzJKg
LfaGwNHqM0XIcetP3O+Vc7A78RHgBGtya2dkOCsTVE9hpOK2f9y7DRM7/my/Lk35
07Vl3/ibZPG7j4o0xOUQezeYmtDPCJRTl0aTGGSBnl/1GoupSvIy4zS/pHUHs59R
GYXODCN7OBLVtjA8jW1B7G2sCUfR3DTyFYfaZftA3MoYKFrTBJk+N/Lbq7CwHb66
WQovX5WE32zZFhwZZ2G26lKFAX0NKcNP6gurcPS/yzj0hvr3Fz1abvbViclndSKi
NF3TtY4SrWnZbVSc1gpe5rRPSHppfgDBSW0l8Pox0VxDDgT9f52qLnRsVNYw6DQi
SJGk3uUt0mKQ8epcH0B0GFlgTYyJlXfHaLqyFTCD7mJk4x7cYC/SkOIZnk+NZ9op
DtuDvJtOcrTx4zsk2meeYNQq+UZhnEa+IvIiGvUzvzP5K6zH7igjAOOuUQDRUFB1
5akSZM4zDm7Te3zsJ83A20ZfAZ79TSqIhn0s1gOfo6sNS67ruvmOWn/7JcGkQLk0
l1WIDy5RpWtMj/ci9WbLiH048vekXKHZQmTLsH/vSLFHfo2mPdZtMiwdnHSAbdcv
wiLk4NvQNC8a6/kIq4caMq7De8MUaS6g3RSrKcClDcmB7bU5HT/IY+WubEuLHCZy
Rjlqj9YkVlyBbCD5QaVgqwe1hEvyOMmQvF7DzkPvMduoz+MtQoYJTEhIj0T0uJpS
P4WBVlIr+t/bo/bWVGik1gjMJdG4SaQ5AqE1aDKxswfZrF8KjW8dNF+KEDF3xDSr
cb6GXw2W2/6Gbi481ax69kFZ1xNXnFDdZKJGtKaI40PZ8VrpF6mfyJo7cmNRiGUG
gaFqSORJQd2H9ROxz13Ba9SZfraqe3eiJGDk3lZADD6l8VzhVQW0G/xVqzQAHoCv
a8eWKERZwS0awy03x/4bD5BnCuXDkmYQsHWSbfhbMTuEjjjqlcQ6fjg4lLE5sRX2
nX9EQIiXb8T886+n2ziDaQOUvsQ3WwU0WcxvlLWtN4BXQuaetkqHzuadjjWerelG
fw2yTwwCp4CM65OrmOU02fDvG50gSxWRVgtPsYZ5ifnBIZgmKvDv0u6haIuxmqd3
fkiCkAxyAaKk8kguW6nCSGxNFBI5XUDATjer+wvqk/QyaNc+3WZFx7Om+VcSxIPh
gQ3wnzpjz0j2MV2ta/Wl2MsU9utV5bdDfu8Y1EtyLHC2ciG3DwQRf8C1yHUK1PeQ
zg11pBRJsMz/krSnvDizF46qhR3pWlv/wYIbXvl+VaaUgf5xmnkOuAXEw8N8N7Ei
C26sOivF7073MMooDAuvq0kBDqm1Li3HhaOrLS2kpjC4+BDMzsba7sc0O67WWidG
N7V1RBqG8OKO2LZ9kEpFAxldFwHl7OdlgMoJuie0FUbclNPABxq6Nc5x4i1BEVXf
IHw+hn78Twc9Ma4c8Hx1ahgd6rDaubg2ebY+V+oe1OzdUZPQE5yTCF/Be7KIPD70
JgBa/48IYPPc9JUI7L4FCW2eCUyYueXU9/U4+Ba/7k/Pa+7lRtCABUSar7V+4CyZ
jTAYLA6wkNgnsdSDOz6/JYTI1cVAfnYhM5RevDWLbrX1TveWTFF5xo7WztqCuOFz
FXn3KtmGDMEmjoHAotcS+zQcNXMfO1ol3oHRBkuIw8FbKR16W2c0f6wK/FS0HTH1
878L5vYPsu30kRdgQaR2JpjUCLGc5mI3eaqMvw7/5LYAlWOzeVUSyOOZnaSnihvr
1+rOOoYe3nRj+0O44rHSwdr9KgO8EYue1Lcr5e9GYIYTtBJnDcFdCqes+4CGMP+z
8wbYkFEJPDFPbKmEygzVCLlOHR7VS4IrUEs7wlvgm0hQdlXDnTSSp24M6gQQwlb6
a1jCMRdZ/0B7QFxXsMQDXpR08uN+ZuXjaDb1WR+GRK/ru2AAKM8lmy7NpUbzC1Y4
VDhx+T+YW7/Nu8IOG6oG3pRTdvnp7hWiXsX04d6X2URDzkEIrUENWBccnIYSzasF
tEmmMDKUBfb4JGr3FiWzeC6XQxRbuueUFzrbcZzOLeWn8OcCYoe3o8lH11evC+xB
C886Tscml77gkYeMfj7QWuQXiDAusxJbfFUCDdubL9PQsx8i8Ltni2YTylaIpZB8
9e2OHxpv1p9TL8DfvspiXj/sIe8b79T/utsIyR+8duqKwFnnB8n6StnBfXMFalNw
Zu+t/YLFAhAy9+tKfman0kiKHf+DA+3viG0LnQAwO1XjEAHW78PSnVTC+hKMyGTo
n6VDHHkUK/IjwBRMB0w1JEZZ3W3TuX+SIUdWHVB2wDbEC4zgwjQLQ9qIoPNua8pG
qnmVMBfq6URl5eHPvS/4XB89x90YYQiw4CwjZQr2rQRdlWG20WJm+N1RGFaUXy8N
G3fmYc3uDkZa8Pw75hY1QMLgR5BGhe/FEvxuxf/Ss/EsPm1DAArHvad5Bjz92IzI
CnutH3H9GjReU2qsi26jdUSh84Ki0Us/GzGFUXeFEJHGM7vpe4JVZHcH0nbzBRsr
rla+qgNW5WLVcnBn7qUBCAXSQzjoJNBy3mGzz6faTZ/iO9O0ruXySLKPOeuGXjE8
W6fTETA8Lz25qONiw4ZTXxCzNR10SM2JXGpKLA3+d8WHreT9VffGkwyVe2JtlqS9
xptCSqiwmSP3JY294Kj+9Y8PaMC8qzSAKSAA91jlGtu6YZoVIXMO1kamPcJICPsv
7TcIJtMn1XulOPPrgZB35zMd5bZ5jvjF2689v7SDCxRvru0FCD2n7MfZ8Km1FpDj
1l9dgs2GOOyqpbOmc87UeA8EG9tX3R6WPzIMNCSRRF0yoqrSP8Ia3RUm7RD7GkD5
2uqN5cZbTzqZgsoZSlHYRElNehKvrny88lQlF8XKsFQG2m1c7+Wfwlnor3YNTKJV
b/0NZM+P43ah+Y7Y+GM17Siui1lkwrce1yvKQ5cTKDtOAD7lp/1bzq6Ld0KJe96E
aAXjhL7ykQmM8Ud9LN5MKoFuuZrlhbYgR3nLqVHNqnVxzZe4o4YJBhsE1ePwvyRV
y+msfipRn635B69Zzi3EPpv3uiFpjfGi1GHPbh+Va86LjLvTF14fkEdKDOBWKD85
/MMiPPgQGUncfFQnE66SqA0/nFfvN2LO7I0aCf/oFqWkvG+qQ6Z5qMsl5mzPXBU6
7lTRISB4DQeQwFnp4Xg1sB/ntvAuYrjYz9o4CbaP782zWxWueA7D0Uu7FfRmPhXZ
WvgtrLRFfcBqEG3kHTnN1MB6jl7v5PGJKC+/SYbMCfdNxO3/sCk+fYIPGnpgA5OD
hUXorNcEOXjlZUrVhW5vmsNdNjFv6WAhY7Y+aHrfLKBt+eaBW+nEcnq8PLpHB8IV
mCe9WKUnWiPVUVNM+0BhGF9il+eu+ARTw7mfs4IGimXqFE/YasbxGV2ODuIesntm
AdFAm0UzVce50J/s7N/AicCAtb8XxujBMAhBlWXnxYAh9AyZZEvPr7xAQMko8Pye
V8MaAcbaPtskT+UJ8zu6YwzEfQpDiCrS/Vx8z7Uj1bIiFk++X5qP6l9/8e8Jw9OZ
fVLxTkNk+2o96Hita9kHHNAuBT1q0mzIV7Nsr5Fxsd6Xyaa/YuF23ErEJXcCkqgd
C3mvgmUqng/fCY2OwbWLjiUP6levb7IfsQgkMoej3A57mosx3wX2es5coGZEJ/MS
4AMJgc/HtzUgaLjzyOJ5dhbO4Ya4Zs4cXpBf8J0+rptiNpc098sCK7pBOiSfGbJf
KyfQmDkNbCBQX9sLtFvybSRkoHu7wWZpU5s10a9sKKmNnCFr6OAGCmKrxTG52lLq
zcEAVETCxlzvFZzJTKUWaQVC56OMBpVgmhY63RGYqQU5OLVW/NOy/KYVc/eP676Z
r4FJtcYTnpVsP9mAAnujkvUIm4BQPZk1rPUP3iqN3nYdvzseKZMvJNMX83ojn4SY
i/YrZiAUBBXsKrEh0zXFNbF2ZZHz4Q/f2a3pS2kdNQ4e2M4eK5Lgqcr677Ys22Qn
yLZBAg5HOrPPinC4AoOD4JD7o60yMN/Xi848vwne/Udgv7SdU5Qn/WaNyN/dO2HL
FiUd7JzeX3DdlmhlY7uCY7tnkTZ10d3dQEnHeULGMXTIQcuUUCWh61NR8bxGw6Vq
dPE+2IVYtTnwu//eH+UXGxwMcQ+ucploPxcgaPeotuvQXrjnwj7kmZIn+C6cPwEF
ul0hIZBt4DtR5XmCSHPkKCjz9Ipg0c2bw9aRDPAbk9c7gAZEZSjAld2DHSPM79AR
h7dwbnLXAmdcnHEw74RSgRyIGv77RKUlVB0AU4zlKHWqhgZzzpPhOnlZ0zQMUAWt
qa2sQMbL99yHV4W7k98Rn4w4SUsXJKTPZvOSBlOjpisovjsU3bxGK0z87HO0d9lp
IhZh4Aps2FryjxF456Ycnvr4Mf2GUoWJ43rxdR3f+SdYvof4fUsb8kVvsuzEvSOO
chCMnTOk3oHhx8z+O/OD2zj7ocVCyVgs99Ex7EUkEZl/SkbfiFBiexZVA+aPJYCX
rXB7Jvs5nojNM3m2Bey+Xx/7osYtKxYLiArcgGHvbbcrLTdW4GdjQZWhidyj2mRv
tL8mx/UuAKWh6K9WevRrNIo+XEZ+AnB1/j2hx84wt346KLH72Ct1982qVoQ4kJyV
Y1A2ArOoD4/7tiZtnJ6LWc/J4FJjfTqIT4K0DxJ1nz8szJLDOEV13TqV9yL5zbZ9
O2DBuW0qBIr7lZHMkX1UQCaXGAKuGAPrpc9pDT702bprffggnT5mYm7tcaw5Mqev
7XMk6Z/rfmVBl+eeYeh0iELhmp5FelKXs1O1UgwrVVQYvVZm1JjaFPDZJlMeJJjb
CERJb6cAMurJj+rglfpmpZukdujUOpHRMdXBAhNa8zlMaCoRbnFc79XEu9g25tF+
x5rRUD5xCM3qPFm2qDR1f6Grca8p9/o/BsBoO0XcqqefzmWYOYYn/8T8SCI8wFiB
QrOxu90lU4s7ji24LHhqxydv3mRtIKH3qniWlkGmtldswO7sS8rrZOuVvRgiLTHg
Ac36MHL7EGwHecryGD4UfuLTj7G/+bI8ZEt/6mWpU5Xm9x3IyiPg85Vq7Fb4lWHW
44xdWv5stbZVA8IkgBvfM1yiPixTzIAUNpmSsBOLRoxCwIRJ4CsFnnYkq8yb9NXX
CnUMIkC3j34MWE0W/PBB8WUe9dMoVkPqBQGYapBqesVT0m9LqeFc9G2rE0azUp6a
wJpCucqRd4uptXtEbR3Qi06SHI3KRtDmYoGVqeZoj60aJXw1gOCETXYcD+PzSPdA
FsnzN0nL2xanhNrWwj/vKrrRlwhnhP+2uFybbhrhKdymuYM3KNkzWln0ajx+gw4M
EtSarKgBMk3jRX+gW9WTFxHEIb2biLp4lUrWC1wluGn1/6Fki6RoR5/tck4Wtjeb
ZMlEe2zbXHtUgNDs+0sEzlTuODXZCnahvI9AGCgEcaDZ1TDbbqnu9IM2wN9295YY
+kSrTyfd1kMLQLg+qW7m+Gmd6WsxUo3UI1Mgh+CuJDoZFVF1mT5osHv9ZHDSYNsF
tUFqz420uFNsICkU8Db/r4zOZklSYVSALkqlz5PC3vBHQDF1zFr2OiK3p51CzH47
xDXv+q3rXE4T/hbU32Y91eJXUX2bSfBEuYPJM5+KM7qJvxwTu9ffuuNVBEeG+kQL
biHxxDpTIj49zIgsmjaysxQimqBB4A0Sitw5q4/GEQe0fMbSpjX8uFEDwt+Zva/t
WDFC0TB64wY65A1UUKY2Sip/9Y+zjUVUAToO1IKAV3ceWrFrhgzmd/vrq3z0LDB6
VWwAiyH/dnC8T10TjvKyI8WlBecz4g6G09GlXDeS+f8TFp127q675fdslnHgvhao
2ol387/aEzmf5ilVU1nx+xtxkfN4hadw7FKr4bKEpN/Lkr+yjo7yBGk90AgikQ9O
qGTzPz8TLM7H43bGBIuVmlmSiURx7ArSN3QhBO1Wh++MPN0INeLpOU8xDQsTIrR2
AHPT0+oFM+XNvyQ7yP0J7AwDlPCSacR4rT6hLCrMWYFRzP1cWPzYsD/gOWuIxg8G
X5C0zbSWGHZ8vLi89OeLvJ8zGAvQTWe0lVE+AcSuqn9SGF0r7rCwdtKNkbL5AkCW
ZvsAQz93bH40X1S8SSn/SZF7mAEUh2KYH96ph4oS9GXXQvkwWvTEktFfafjFi0aV
jqUsrHXUjY9GrhVg3ZLNrKkcvNqtjve817eWrbyziOxzncAxJbJLMhuHgb9osuzA
ksrf0vwBxGKjap/mZSxp1EqTi5icjLry2cr9xFSJn+jm5uTEYBrkq/fBp0BRyogv
7D3fU4vLap9uyct6H7BNchN3elRSIRRy5CfHR1P5RHaBnAMuTxLL96W9nCwND3Qr
E9een035Kv2EwRmUy8dEUY56G9fKVyUbwqr8Rz+k6B4U8Chx8KK3KWz+qFkpmLI0
Vy+RMcz1WJW0QftF1BrxtuoBS9XoKAyZ1aMgiJJYb4n9oCh0LjokZVdXzJB5w5Oy
7RfS0CIah5xTFzNrRc+RA0cCyd+qlE2zdBSyXLGXw6ZkSkrUfkvROztEQZ9o3PSd
A+Sdk/ZO+G9ePbcWuxjFGeLAfIpB/ohqXt3X60CzmMduRVAjMwo5PrevZvMZlTVl
QIJqKY+E58YDwZTQnGq0OZ7s3ij2OaMEOTmXEHA0LoI3y90B+HNFG7PjyzCI7WQD
JvTL7GBbEJBalsx2tWj7oLCra76t608+BTRAHWjWHe95W0Ari6QL97hLufPE3O06
TVAh6pPlqOYTAtkxXgmtzlRjyMT/3tOE1zSqrfBWIY6B+RkGQLmuoeRy4KVeCpiQ
VD7LEiYPGQXP5PofVcodbL/vr8w+yEwIFbwbeMlGdcZH5qIW72HIXI/wvVNPxPpm
Dz7UuXpBVtV+deUDolNYHCV7ctaJdD+oT5mEjCdQdHA1dkaeBCBejz+H0PcMMBbk
ooDbLp3Si1/IQdBGbhcjf6mOEIJsdyVdoBJxDqiR43RDppypdh9Me8SRcEys+5Gp
cu0njxYFloaSs/voayPc2opaKdNEp+35sL2erULezTKFZsRhO+hyY8PT0T0td1Wv
dktf25giT7IAFwiM3O/VEs9zKjAxQoMUUpzxIrhWFPf4bmEOLeqtFiZpF0v1BGu3
camwDRRVZvhgn/Wr6wa4bDcBFUL6uk1VwItTCKYWvlvQVDKMG8ierpqrPhMUTfdX
eBc8mYZR6m1ok0EbA+CmkQlb7QVllNvcGOnaFv9P1uFdTEO/2R6M06/m2FK6njsd
Ra3vL/zYW2unXK71qVJm1Dtbyi5Xsd64yDPTWLmj2rv7HdSBp4rk0/J580Me/pWe
TidxUWLBqmV7AuF0ORgUzU+uEalcqxonPtK1n3gPQS+dOE1HSp7aNXVGlFBquyw4
jMhbrENK3TtOjnDKB1HrK/Zi6y7hKA1P1oOM4aXzhSGAxQQLvSTPS7jkKk/a9hhM
8uq9rdvukiQzoDYCaIuUPMaSOL4RxOVW8lHaN1AC2Bc3K5ncVqZ9oqo7qMJvguIp
TCHn69eKWMkIv+jba3y45OSIxLDU/9kwYDErutdvhN/Z4DfxxiF4MSqe+n1Vy2zU
8ZuKHx0qF1pxKMr2r5CLOePFeGGnenNWMsfKfBby0F1rJNfKQAF8BJzJM8JFcOSL
OjCdKmDJjBh7wMGauUISGwdOGVrugd8YZUxOlcI8v/ywBHCnSOzb8A/vZZLfAKFy
+c4r+y1P3dUwn/GYxWBfQT+7GUMmNXjmKhFKWbHJH7pgveW4V35GejN1WFn5Fcnn
w9Yvhq41078L+3sbtFvZdhmerKpp1uy3J7PpdUnAPhbDi2C06IkWt2d6haB1iUJW
qh+KnFJndUYsyWw+S23w0ZnwjE1vbWyvN2ynbouHtEQhqfQcJiv1ecauclBB7mDi
chSL1l0R4y2c9bUHdtywJLbg6jwljRRIouOPlDCi0aUqKm62SmlAhOYIrIAZ3Kmg
RCq83Yb7ybEATmHL+Lzkq6wJTpJf1+Bi5V79syAGyY4NJ2Yoo1VNda3sRK9QiVtW
GGcJa38HtNY/ZLuG0JUcpvcepBRi/Dtv+/18DI09ccGdnsCl3ZnD0f/zI67LrdPG
osLrvFQHoiSgESbSyHBiWqr2kxI11cpZnQN/l+LbamH82qYfbDpc3GCQuoOFRJF5
JbhWW3/ixFcVGB0gROrDoqnrMenHPBf8jymN8wG9TYJ4s7vLurNm53iYwRJQ97Zm
fGbFQcZY6g+3/yp6qNH5Muc2mHVSJz0jfE/kGDyVWyjGfLBY1+CnZZz16dN/Ibeu
1s5vUYKXwb3ZbI1ozr0Uyqt2IC8SVbhyaRZHkQqo9pVHwMSdax3cf3nkm3mHGmQB
YfsnWNxt/TA1abBI3QIpdhqdDF56xGUJ1vrzV2oFJxFSscr+0lWLWgvBWEaQnuB4
CoIHU1IqdLb8y1IYvY7rrwNmjljzZI2kZaO9D+VF3CJuzorg74ljRkCyTEyZZMc1
gSNPZRTvatslySgrk7rGIXmIbCby+LtaF8iQE/is2qhPQTc692ZgbbOQcT8TGmYn
`protect END_PROTECTED
