`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HFoDM+tm0l9FZN1OVfrlx8DDPdqEbRxsH3KPT3jvfI3RrU0k5Clkh/FfxxZAI9Du
cTJoEsgM7M9nrIt9dj97BAGdjsx1CA//EjUmLALgvg1x52rjU5eDgJL/GXuk5b1n
gRjKE1iw4leS7rQvDCvue7dV7u59Mm2eG9c4Yhz+sL7tQ9dUQYUfIZ6Lt7DkJBc0
W+dLmfZJPd0xr5VSma0GsywgDqxEvsSE3TVHXD+KRhXvl9gQqzQ8TKa1z+K7QzNw
YNnMmlNGF/jfRdojq2OKTO3JD9/lhAB1dMrpnlEr9UgdmuoIc+dDHNzQwcY1y+HH
CB3IPkxC+E2IKw4fLCKjzqeAU6SA/bHMPGQ0L81PucBxyvnWHzgpn6cURup8C1SO
Fd/671Sa2rRMKzo4rJmbPwUaNh9qhAtMN1HJWSWxxOEu5LmP9/+OwWmRuBrgz5lt
pzGKEEfQouPzhc/I7MPQkTTThUErizDzbqLHrLVZtLgV9EqipnaOP/fq7AncS1EE
J0caileArx6PMBAfqNu6ljem/pqr1dRZexaBuIhxhdiK4Gyw3G+JjV5NVZFf+qb0
kHdQtoHoWjzsL/zv4sUJlhzZK7I4+DAD1f4E5PmrKXWx3bpjRiyLK31/1/rZG/D/
eifMv4QlL2ya8qt2nHUhK6daFamFuxI3CLaCHpa4JPpbXWB/u7JgFM+2poPJuGhj
i2DkAgtavrsTbujsIhMBOYI+OFFxHLxfgJbIp3WqCe/KpXx/cZGD5voLY/jfc1R4
0Nieq5i8tItRlD/p/V4xpmTuw5mix/8fl1KYAyFWpiwKnoCw3GLp18GYmnwDaWM1
bHx+SxHTLxyOm6yp6U4rBE5QmlYwFcO4KR7BLPMVctZzVM43c0Wyi+ErkTMVbEZ7
mJ13RYB6cFq7vCCMZ5QZ6Q0Ysdn+KsNaoXzs3Q8+Pjfe4Wl85UutczaTF0cHeh1x
/4jTJA1Cl+qvXWOH8fWcige5rU/qIv3QAFDf9Nov7TFbWziEw36OZmWcef/yfjE1
52e4fUjhPHbeYr29wak2xvpcAJhJ7fvg8G92oOUGy0Y8XCOuG1sKyr1CnFtbP1CY
fNZ/zUt5WOctABRi3V9tWja2eskfKyC0e9mxQ7wrSo/hp+0F0s+hYCoPiHuDKrPi
ehMxUFIzUF/X4zNOKH0qtquJVHBtz9Ws3j0OdhqdLnlOCa8Hrq31O+E1uI5ExdW9
fGwFthMAHS1wBe6jD975nysnb1PE2Y01RS1UA6jpBmE6NJmNssxDRJZ9URuuvcrC
ChCbm35LiQBJAnr1/9V5zSXz4dVKuf6p7s9Yqy1W5/BUjuSi+kG5gM7KOLP9+LGB
e9YwzY8F+zoBRNYuwvBU0MN0Jf4DUbCckEsN1iPCwo0oVSEOi/4WVzxLDUZeoj56
6tmfAZWMX7dFaf7iJhLDUw2tX/Sg54hgMuUtWaNEz5ar6LCEFzGFaU54Gai/LQ+2
YVXSH94nTxBubmbTb3QHJU9tVY0TYS5IZniDBm0VS2/ocUDsiRp8bPr+WfwnG5Ix
qs3EwtueXNIpqnn8W/djurRsUALdG6DIrP7lU7VFvMfdbyW0Z1GBhOgU7euznLqz
u3XkWAhaP5Tse8w63tqE1pora7d/UqS1k3KpNz8Kbj4E2y9x5oSTufVkzchjZ5zt
zXQOTm2J/P7I9c5wLkdT6usjj0WTkukkddlrJsJXpnwKb9maQEp6MjO2j5eJS/fm
is3V5xgnrBw0YXfdC1TgBspJhH5hbLlooKrx14iOFsjgVA6LAfCIdNvQX6NgZamD
Qw7PP2fHjk2gi/LYWgahWbypX5Dnq5nWKbRx7kScvo079WRLXXeCRKPNM+SR1a2d
MoQomELn2KulmNM7npuT17vagiIfLyaLsacK8Yy7FaKPsstERoV1SIcTdaRC59yE
U0rEkO5SGPZhMbl4XP7dZykn/oOqAuq+mempMqh25VKX9Ft4Cpa4TFY8c8rZVWJj
2QeeHSDhwXQ8M6rTan6SXNoZ0CUKu3uQ0Vfgr17PRXvV3QTTEMdPk786P1N6NI9q
812lIm0U3SiJ2tAOhTKWy5pzQNEOEwdNY6ilcvefE3bIYupsQn8KgHr3MemZpllj
fWLD14G5G27GyuTDiS53KgfZzWPEdc8KjfoUsnKYnbPZD9inm5ZXngGC8Wr6e1YL
l20iHDdzyuJEliUeF7LAQdApTP/eyR75D6rKLkUquSYfFnfnJOVhvsI+RFMNtoNW
vlKO9oM1AEeEPdvyxGLnthUkDZSHVd3yxcCkzgo0bAgVMobGXzqVSfj5I5CRK251
dNjV7AtX4K7ukjNjtFLMoinXCKGQaOA1pIgvpaGy0WUgf13AUDEEXFC0qyBCUh0l
mvqolvdcerhFvQf+UQXpSAikiwSNNhNaulvpdqSWa70w5eXa4LjsXf35tOWgJlIk
fzCoiboCwatDXsHn4yHA7hFV9K6EWJ4OuEPaqSc9cufdHXPSW24zj0wNSwkSBvvE
Cx9s5GFSWStLAboZWznouIunYfn/x+WcqNN4eRTMnCX0lNdaSAf7idR16VJEVL6z
+mhzyVSDRbTqhPeoeVhBlrHfxTIWMD8noqvwDwA5O9U8m6aIuqLgs9hcwC+jqnT3
MdMaUhTDwlr4Mwj9kfnd1puSL4n9R63qZ0ktyVwsPAose9fi+s2U0xvC9JSEMcpC
aSmZRThYijfnHxFRwQ8np5iksE3PDnmuVsTzg7w/zRQ7jPyeP5ydkpWRYIX65wVJ
MZLH1HoYPReqVBxQ/vvhrWHtOqZ4ugc5RYus4/ffNJ1FGbalQThLrNOXk6XMjOAM
iKo9xkvteDbVvLnF2EgToMmNsxsFhZW5l9rn9UYw6sJueDv+/qPfQOQUzHg8WBwn
i4fNGWXOxjO0lzo52BoPhMLcT7rzMgax/6f2th+J0+G1wCq6iilaP7pddR5z3hGC
fUD/UcJL6CGKJ7zelwzytl4XbTLXvVbdGGqwQ0ZGYVGszCULzB3nlcsx4dIoIoq/
rOPJ29BjUR90lm35ROHuYvchHgY62La/DO60KuQKFW9bMFhM62jxBtsDomLxIpRy
bxaByg209Am6AqRrTUg/YVgnga8nlvDRhX9uXguF+m9yeFTrgA3mwR+5GmnCbk8D
ZaRDT9otNX1Sy9GFKKA3/pzv1wssCVX8FUcqtJq8S9oHLUf+BKY3cHKU7/kp+F6+
2wmH4GPHBGAvgF/gAbY6AiOc7Z7xrfBGNfeMcpgGxry+S3WhR1GXU6mvbukwan01
iNJd1QEoyfcde7fJ+nTOv+HDJMpWRNcJJcUFUR0xHwJ7lDjdqr1s3wXdaQfFEwWX
3FB+zQabn3tbIl/ZFaMEDlqg6QCJI82mOKA0/GoDIvd40vQ/hzdB2EgrO1F8iJfw
ZecIgpJt8xfZE1bua1gEe6ZSv3ygyuANasB7sKzEkPZqXFVRwRN4PPwBQhaRZSvM
RR7AbMwvnzt3uh1yrVLu35XOEHjhQ9wDXVRUxhh/RRpbGJwUUkfuuOkocyhVHThj
jCWpYfrMm34V2UOxX+wDfXJ9frDTRA5d1sWY9NdfTdzM0m2oR1G8WOliqezvrIfY
QcseYVYAtm3Lod185fjm4i7YaLGMhFi4NJ6SitZ9E3w9uO9HApBPEaUiEd8vpaOE
95AdvvUlblidXiZz+BUGc0URCBJErt/zOFjiZ9S8LzdQ/T8AhbMCZg449usr84XE
yOeuBqrs2g/ieXecX8BZOLT5uGnpvSd7vxJ/mQDRLBGjTQEusR46S7WzqeWLd0xO
Pxprg/OxD7vXBYOQCaCTDIsE/zRlCHi9P+3gwn9JKhgEUDS+PwLXvQbcMyxgjhbw
kRPV5W+I0Lf3aDyCT1kqj5Sh8DC0MqqVxNNdvzosuUNHxUQ2fQkXZlA8YTg0oR06
tX4H6HHBrdW2anUOnvV0XghqZPFF4IHqVBohoNmLAQaaal47rrWyeE3R1EAyIYHu
YhDLJA0ofHyM+nAXWc/t47kY5EMswLLy65RXCy1+xgVvtu7Xiz+ugbfcqFkCI4Cn
ziMTF0bOSftA78qBEIYlMMY59IFXrJxENiiaoyYEa6qcw196KlOu0xb0ouc+n1hV
Wfa8jEhI/PljUCCdBrZeVDQ5Q1sJYF7HGuAanK8PaRRR0p/xx/VlELomLts5AIXq
vRskPFgx6WDGPtrV9TMbmkcg274vd8fQ8w6cQ6h7y3LezsI3JY+gQFlgCH5ooKQ7
dkgIzZEb5cMdIYXX9HYG92i9dB6sqruI+HNkNxR1O+bP5zQOejyrt/SbUicANvOg
rry1UusRygMxkK0+05wuRxVy54mhQCZhcvZS2mrjzkPuz/GhbWsspzPdp3pYHCtw
1BFgNkyfqLmV0H8so6nuR1LgaivUlokRR6LtfJe3FMGE07MLAnEaagzdc2b+qM60
A/mgleFi1iYs13mUaWloEU8D73u3OUMbHqbt5RBRRRVuq2lWJ4i19Nfr+zr+a2jS
qeyTlhcBAxl1VBhbbH700TwpRLiu0jP48gbqV0jux3UHDf397OqoLBdxYyPECcM4
EmiYUarBL/FGTL7mVYXWTRo8xTDLQ2jVKJBE7g8go0W+LbkqX6jDNfxyjnQuqMO9
8AXik4ec7aEmjww5pM+SZM//vuFgMpGNmiE0SqrbHLZ/W4QiPOEuhhEmxOrsgV/u
mPccZpXtS6y8YDbebl9TkHW/JMFMOXnzlHiVZ0Dt4b5rropIA9ztQOUJo7NWECkm
wOHwAIymerB5thF8WpsfS7blE070Gug4VhVn4YxmDQPZUAuO58Gq4WYjwGzxAJeK
V9XxxA4EdDmlxgGwtr7nAjnzDeLmSdiI0OG7hyyoC2Evx2q1nfulYXN5yPUaqE7Q
XaiEXzmi3onf42yCA8TCj5rF/JU3crOJvmOlvvG6KaeGFtscznhbbLq+PZKbkhTU
id6/qQehS+CFmY0+8VRDWHfIDsZaZfDeibPkkmMYYMM1M95w9wa5yeuORKejLS15
hvjlS1x4lsYCiBWuJO09JcHqe7MJjjMQ6IMeyCnLscrx7s5BpZ3rFdUoFiPdJPni
n//hi1W9+l4ug79K8vhpCMb0T+wb7edYMBkG2dJIx9rxSLzsIeIj8HW41IKSaXPr
/jlR1EecrWiDKV2TEjvz3tyIor6fa8gSe1OOf3B261/llqa/0FXorotuCyZLz5u6
d/vdNc6nY9dt4eKyxToiB6pzOQmNLthqdF6jnYuYfriveWd7WxinaXjWH2OJ906w
5YnqMnG2RTxhiuzYiIuLmKKllsX/nFe5O4dC+TAPz2Kk5af5oSCSliHn26WqiT4r
lECfUF3wPGOnikqIZ+Yyd9kaVQGxMdcWRdXs/wWYZrLUojUXX9xv3EG9FOv3S0yv
elv+r8Hpr+TbM1OwO7zCgxZa4a2ZAHYKahQ6HTTHZuRNhhsoH+IrrRqcanSNWPUh
YrTRLSFCs2pVCSZznhZ2le6XLYAKlEieLBxr+3C4xZHs5EWv84Fxp+nsCF3GszmX
RQ5W4tpUIZ66i5c5zyJTz3Op9zUdVobDGwlHy2FavEU5GXBog2eP5kxW7I58Qipl
55rOzlKJHg4UatVZMe5A8IBAGsPWw9DHpeXXA+Jo5SMgUjwhTwei7/nwRAmarDAV
ibeMgijuZwbaAeHjnVP5yKPZhrQK4J2hGROL9fpazvbuZ8w6x5hMTANURa9lzD0h
KLVyKM3H9GPYssR4mgTD34b1J0Xiuc4i2d3S1zFZdHJuulS8yuPs2jvOdTFh3uaA
HYizt5Ao5stUU4vpkFHZE92kymE5jGOWmdTYUF/mGEjYADFRp1m7yI227UdSTkDj
Q2UU/hNhsl91hrzntkRSqTaGLT3cKY5jpnlRc75BBfsxD19uQHJ2xpK4vOoWFvZ8
UnLrLioydIDfO9nwgQXg+51uGrR559CMAiZR0pH7tjljZMctgx3VIbI4yk2dXJa9
FlEUt0EYGcABV1ZL+nISqkaerPCt4NWXvBXKQnqADa/8pTc/GeGBxYnUXo0p5Q9q
4EQDxGHZtMDxlgVq2AORRyWntZEtT7UJ4hlaD/HZiS5Jq/At9wk6SQO0DCOp+QYZ
iufAkR9yay8e6RmHN5DqjLOFkqxUOrQD8CFopjd6kLZhzhllTpHYEXMDS07Dh1TJ
IIFTeJaLdNm+ih5aUC2fSsAXgXKTDMFh42keSA9uJhEgdwZLpCe1S3x2Ymb2crnx
b7DiAJLUa1HGnTaiasRAt7l4G90nUyK4ixQ/Z754eI/z3+Zj/7Of0SKGWRAdFP7X
8+P0AlL0GdDnLOzfRrDf61H4tzZeAxsoeIHB3HmxanF7JUswLPkbSjCG6BMvNQ6G
PYZwruWGbxtHX591yFQwtCpJMl7mtWH83jUiNbydNApRshdsRmdG6vEldiph1C+X
FtdlsvF74d//1i5/UsMF3NdEjieNSsqe3e89/dQAE3gBbk1So5XJBnxhHvYrt9Wy
Q4OEmR/2ZFK5J6NcQLYs3rsKlq5aGdk88oAPnv5AW7i+G7GNJk8lxs7A48Mbzyph
BGoJQBD8P9TH2hAofFeyZl6pKOsmb1a/5TxPHy864vWHYxXdavQngpqz0eFy+zVp
GuJCz3i9Vi36boqg3ehbUKF8KGh1+Ua7y1d67ARLCLdstah1iGKLXHJousmBgwtD
bHcUAw/YY1hfB7UPpR/r/uNIo+chTfkiTgbFCkikQTiamnO0JE6B2IFdWNh7KiCv
VcVIGz2+k29aQw0eFpGBkh5vaWY7XaJlWvYQnqpgilwe7VSyXRj8Ptn62l0Bg4KI
HBwP8pOnDTEc//MKreEh3k4ZFBBDmFK4BEF1F+MH8oCTyImqtTC4Q04I64Uyh+M9
bZtq4eg6p2wjoMXEYFiLTBQCw/My9Dr9qH/VKUymjWkhx6mDck1WP9wKu9PVgk/Y
+fkQWaFZO8m5rn8wkUBkHp0gva2ppKo+hYI6W8iyiMfsZrt5NImDoJdEJliY+q8d
4um7O7wlAICzuU4SRKUhVrEuuThcPTH3yr1moAuZErij3EV47/niOWmInx4tR8VU
DZroo7VGJmIjy5WFhXN3Hj1PBdIZNibtsGXeTIm0HMGvgTgIPwfxFJucc7/xUBw2
Sbaz8c2/Noa43ajBGtYcTkX5Cq6CUAkSsjzWmCStoHnCqA1KO1B2Nm7idH+Q9xBd
0THukuaBQUEZOK8oI9oOVnyaoG84iAq4dK2TK3XlTCvqca6EqcD3OCgm7oJxIBG1
9wXxTRQ8jl55P47ztxp5YusWZQqWC3PxIcfx8opLFuSU7tRVgQj3EDdzqVP5L8+y
+oCETn7VRtSmzx4hvzHn9WfKBehEdNgIsiDl04pMmPXE54zozZXHUjNrlvHNYv6P
v0GeiNFVZa6bacC8IczQamT1ORrOXZDLBkEP1wl4hKHso9NIYSgNTsmAeXEo6JV2
a7+07q7Yb6tklkZuwhBxgT51gSUtQf0MiKzO5nZdnli+l4YSjw0/QlFuhoZwMHdB
HLLmDo39SzkFheUVrV76ulx/vprwlWkg6u4G7Bl29AO6s++gYK/Xgum6Y/QwZ1a6
wmRUr4A8b7+/L3n3IRbCnnWpWBbSatWPOZY6YCNvCvxhU0nMwXA4ROmihB9pkEWQ
KWIiGXOR70GfTZ+kidoiC0C/cxjkwp3yHIYE+IEbzZoIBHGPNCLAPWUqwQAoaqVx
IS3qVHqDOGost9PmKt0/EFHz6wuXAL/uJRt9B/2t5NeKiu2Tlj/Ey/34LC3drXBe
RCiCXM8mq7EFdwDK9IZ30hhyyWKKW/bGwPtUM86uTuGotHimglc3NrSYN3SpNBiP
C/tNTIYMmoY5Z9NuKDZmBzSjDLHPTgpTjOQMdBIGBNxQxR30T9C9Df86tkccdcN8
UU/Pf8T4VnRNUw6/MXDGWYM/vLYLi4ifZxfO7C1hxh7aXpXn8K3AVFNp6cLoNAVN
fcJIMOKMap9gb/c0tW8JpMAUmGCB0oUoG3UFaIHV3r5lr+gJ3crKjQJr9KNx0+u7
YD2R74rfCVTmr1G7ieh9QPs7GHOAvct7sPKeyKQqNFnDJI0HjQQJlnNVvdDcobtN
j7UYbUpqsT52EsIbEicx6t3j1oZuim0t2RpCDon4D63qfpOyIZeHzL7Vbu5ShJy2
2HmguoC/PHmxdcLLfDRsVSSqawQ6gZO0a+bt9hQMY23sJo0pszrpn2Eg/Hgi4cgl
hiArFLrcKpUEkzoIKc1AK3OzaJ/TJZAS1fh8Q6jUE8ZcR2okk4pYMeb3UuofZJHM
MnXFZTJAmfE9ayyxZ/+naZpBhyk3MZDlrNcmd3WIMcF38zl0msa5PYvqMquDirEm
Bt+VM8LA/hFvzOJKKIZQLCPW1yoRnhH2V6QYS7+sVVZ0oy2E4OKV2k1NdI4vfTNI
cJCnXe1xPXI3yRoNwBtOrOs9RXlT2MpOb2GmBC6U8t/POzE0iQ3OWvwWallo3Lmb
N53doaXp+NKvp9il+mjehGlMS+hoiRfDNgHG10/N4Si3g5Jpocan5SdUwbfdJqWY
A212aa2w+jP5bUItLXiDAM8FnXvVipmehfE5nnzyh3S+Ii9IRzDZH1Q9zJAQr7p9
J3MXQg7Afjz6NJq7b75K32ZBZAnH6CRj3lNLoCWxvYbPfD8EwojahHtL0k4PeAAD
YDdKonCB3yRJUKRlB00AjgX+xDID18xBD8LsbCQKzwUqxIVM1zqXKu2t50EMwb4Q
w5JuVQgF5dVkY9PKFbCW58+hHiM36kvb0CtJpQsSpU7GX2Cib0KxZQx9viGpVRhq
I/J3xYY7lv5VlqGMA0PUARwzm98RPRs7FElUnovvgMy4XsN4B6kFZENzCiHylcr6
NEWUGAJRA1n83HqUf3gaS49WDUg6wRtX2m1g1H1hJOr0A2B/+3Y7S/akbXS+gRMC
yRHQJwqaBG/KSTmR9GxyxC5TNq+q2TpRb/OY2axUxuwhMS1uWpz3myH7ce0KrF1P
pssOGnr4QwthAudhBLMUefJex3DP+/D5HW2jU/xJYSc3K4+BCzxhfPYV32CHCOCd
qW66InKW9R+E2f2pjci0RS/c5oitHnb05LrXcbCe4se1Lx8AwdnZQNHvibp4TCsO
N0cydnO5AFwmZNlgS+sLs2+XyBbEzBDpg7MnEF1MxaDlxDKSelaBVb6MsDZncM6h
u5Y4zKiKpk/wawWbB3DJrQbOM222YiU20t3zYIxdUpyOh9QQz5N3e239PZhUjQPU
wLgLKmR+uyR66G9vA73DgES/+PHKEjbzEFqF+d7sWKg685lEnNtIaKFJ6V5buLIJ
C57PDTcY+rqFmV6fwOl6jjnKf5ZGORSmGmzUJxASenfksrXV9HY1LMpkrQx4XU7H
gwD2Z4z+L2OGZ0PrOMN0dm+B2zTj1Oeo9dnrBSB0RXB1Y+n/xp099h7/n4u1JB8z
NzPbjn0JnoATQrQQzRVSIIbckG9BKUgeHzWz+i7oEA4qwLdcbhntEVz2WPVD7CC/
QI1veRnOJPlAweg+Dwpa+6tYmSFYvXmdLcsjeXvw1oTKozDR9o19mQ85y773gvQC
F5tCezvmAsiuE3bj9mVzIDpQkXIG7JNqurfJpRxsh4Js43iOqBdnbmVp86LptHfC
CVDEx+W5PE8ymEBfaI0u2nEFx7vU2Z3uLGD8epEY60jf9Jc9U+plFFcImJ6TlXWe
23ZwmyQPuB/K5hmb6Lwf2vRauTIN+FttkKKe19JEheA4adj4XIgYxF+/zUJYc1K5
H9jzXS2cLDuz4ZJf7XWmSxoesy/4dq8aLgQv+BLf9gI45dQPM7rYgRJgfzZTGz8d
rC0mlBB8HDXIzYhlowYFEXCTEiHUgSIh32Vyuvv1A2vLfBJUOuaa0cHFSl1IhwZt
2mBk9nstInXYZzTEuGdk/+fxqObNQ8H3V7AXJUgpvJHietZPXcA6MFbuF8Swff/m
3rjmhZmbdJFYuzrX+3jtg+pL7H3mAuUkGJsB8O9V8Wt5gdFmWhDc2r6TgfgJPjB/
LcxRXgEvE2/9ghHv8V4g+hQfLtaVT8xQj6H+1QrTxNR4yQJClsbui5g73ctO24yi
uwqgfCeR5KhcJ36vd6vQ4SFdKjrxr9q7w8Ad6pARbU7M2TFhaqzMs5duz/fUCZ//
aQnFvgs38qidfcM32uF309LA+XjrpyYyO2wbCD0begExJK9bUgcmAtF4Zge7j/ha
C9Gii+Ggx/y9KE7cIxcqNh+JSGguk6UNgvCsIKm1+jJ1uL1fcPOmZUg4mLzNRXiZ
CLQnKEGuPoe4NJBpKiaZOzUHX/ZndSVc7/znbyVqj4QzRblAMwTOFODqJNui7zX2
`protect END_PROTECTED
