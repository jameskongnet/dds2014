`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0lQcBDTmHe2J2k3JVnpLRMiWMV8W9VT0okBHnyWlRvCUx597E27iywm9q994xSBJ
oXgGpBiqLF54Or6B0nr92zm/n3BuQqDx7bLBUwyTLMivVLH+q3qoyIGIiFQfysDy
HrwRKRL9yiVPAhDGuGqp65+w31J3LEk5Te3zCdfx5tofa6PfBLEx6EuggXX2nZRG
Oehsw3F01Iyi+srXkTyHxocgzKgElP0dk2qr49S+kRrHAcR5zHbQ5r+4i/N9d/tX
7idPV9iY5EzRZzNUKK283w78WLYw04ZJDTU0lIyq4ccz1IMHiFvjBnpm07xNfYLZ
W6ow082vzzb+l8FHSQg4asJjFW+FxazfPypX6IV1rrSB9xIMuip5a2Q3lZPfbiW5
vF53Zq0UqYtMrC8GeQ7eYQp7MX6cGzbab+qRG7O/G1ZbeFkHrgTkMQX/7PNTAJoi
oAes2+yp2HVkqmZvX7qxSQcL/aYaGp4rSV1YUI9xQm7UQ64YuIwjmAUBT317fDkW
DWELA52dV7g8Hpqs4X2eeBxFVcJ/hInf3mPRQw34gD5uwDMIVKaLhbUUzcaJebwc
aHRMePfXqAqn9hPMz2agAlIJGfsnMjX41PXrLL3I9rYSDLC16uic6jtQFLCJYaPM
nCCgvu3k4AC7kAtFj2f9cNyRLA1LyRDboXOdhIUWxPoacdg9pJzeiCRHpj6Mw8GL
Ru7cbtL8093aTN0+nBLQ+bi1G5ipzy2IetUPpmjbALr+2EmeU/1A428K9GgLDCrU
IbG9gf7iKBPV7+io+U2Rs+uK9hP2NeoUuvFMI49zqWoau/nrWcsdaSaQcNYgt94A
`protect END_PROTECTED
