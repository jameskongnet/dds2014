`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zhIYoIxVQOB5AQgfGr0ElA0XsU6vdFNP4yGObcfv2Kl8PudNm4kWGWmeXIvUxykC
WKWA6VxPISxKwZAHSQkmXpTaESs4HbNr9JYdZWSbIJE4NirMoLq5LSC/UbiST0qM
+HvqWwiAmnPH1CCkmCDaJykvAEIJoJLHCaY2e8IRsZm6lPpNmxSj2pVbp9Gzb5hM
pV2p4jOfheoJ09kNp2P9jF3y/nTZh0XLwgKIo91cambja3rfT7Qg+/Cya6ANLeZg
vgyNVg834C3WzY+CBlvVEN+tfEKSc2caIACMXjcrMt67Z4w7jXIWyKOMrSF7N0iw
weFrrfQgym8s1lrWhYRz4SrjTIKkOOs227eDZATyxFwSm7fi/UkNETLZNlNg9p2V
iSYsbZsjhnRhsQ4+iPcrv7fsCiB3mV2mgGylYauRKaeP0AnJ9dpJs7LGgt77Uu/V
1nmcFHddE88ioAkpky5DiA==
`protect END_PROTECTED
