`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PsH0PKQqXU3Lv07EAkb8F/0lc1mGThd1WTDcXRTCrrsRXwADsLE+f/rgjzk9hP0+
LEEuIZPcBTjvjNlcE2Vl9ZZePTNFmKtr8ufkX1ZXGOd7XgyfjXpdzsAmfE3GIeuk
uPRPleIpbt9ndQjjfCGsaYJQrgnMndobPwToVBPHrEKXBVYZepoTPm3Al6XzIXyG
KsXtUoXhJxPRmeLUh6vwyws114q1dGOhl0aAzR6DH/W/PJnvKeNAXfKRGi8nYmGO
2FT5b1ikNaxgoQ1k8LC7j56vaLVoN+CTzJTC40sdfmP8NWhc3JJqiTStRXlm5ZFe
W3rFqqCrKPYA82eKQtO1AXBXt22aVn9IPozJ6WRu6JHkDDcWKnhUI6FKglVJ7pDL
OzLLGIhVgZaepa4ePK5ZdERIdvI1KFUPWOLP375dH9Wm3fkxp77Hz0maZw0W0eOm
4saf3d/7xvziPRN3UKux6tBDl62wS5QrWxsLpRZu5TqdHYvqEge4GW/vVlPoi22R
ytaPo1jnQ6UGpK5diRdhwNhlukewi38b3nshyTixRtgGn2LAnnohiWqJH5BgcJmx
zOCtwZUmVCOaStpk5MRdzOfDWSkJIzgzdohMhk55fpUI46LfoKUIsyvna9624ilz
Tzw7SvhrqPDbfMoJdJE1pkVktOkMzkCfRKLf0RYz33zitI1YZzfTMI2Ji0DrQjcV
OdfT/P8HjaOnxoKT2eTnHqt5DJE63KfQtlnDcsf3nXU=
`protect END_PROTECTED
