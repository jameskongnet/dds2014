`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nWEG4XKAMeP41SxzE/zNEg49xBSuf+VGHo0kl696ecskS/jBPojTa403ap0P/bX1
Xh925bs8sN7rMZLOnNglKAp2hSW1wNAWXepMp9uF6Nhop1O8zTsnmTF63LZMjXnT
0Bw52DrkIp5JcAdCHaqKD60auvT57N4E+/qbQY5UEPtldQDaiyMSPSeYLaYhPpna
nD/HfYn0RhiIkLigunTEQfEyDxX9fgD8C650T3q4m4cBHxhiXVdWDa4VAEPCjm7H
WdNI2u/spQ4yTKxyC2qcsryHdgt7HJ4D9TU8tNf7yN4X7fzUHK9AAlLF62MwsbeY
7HQZZkZ4AoI/Fd2hHlwStog2p/WhbP+dcrG+rXTh2eOQeKzsF4CjXDW00LGb6qUD
BAG46rXaYKhDd3WPSwqJXIuNApqPWs53bPnQEJ1rw8JNU8erI4s1wm43IDUXHNzA
wYsPByNBLDsqiya0waKNqyR02OTvS/S69q11GawCpfCL6diJBzhn8RUPJAr+UgOy
k4gWKrDsCv5kp2/U4QQznNvf8g/fjTXbmd/IMW7FObRiG5R3Kpg9XnCfUAXPjPUv
5V8k5MsaIPXHV6KS3b9CMmHkSkUmZ6xPvr4RyiCZvRiCHyU4jtAtlEGb2Nd8xm7A
kABo7Qj1aVQ7C2h2CBaxZNUP746Owp9okaKFMc4c6dW1B/YGNANq8b4oXLD6kbDJ
8qouNHsSn6tGNZQ01GcVdQfS0/4OCo4pJJly/vvZFiY=
`protect END_PROTECTED
