`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GJ8MAKUbSZTaH9XPXZBCo7wQcJZmw1NF9CvafVaTh/sE3SJMezzxaFxB3tKMX0xK
n+OrGrKq437QVkymCzb6tVjzRVB+y13D4bTSIOFZ/wbOg2uRJxv8VWCK+bus17ND
9Ni7A+6LYW/Ken+nChYGshrYGZHEMTcWHOyLD3PxfBYtv8tRkZZG83upnyyu+3T3
qYzwSLfaIMMVQA3tS+H7W/ySm7IgW+tpK8ppOKsVep9idgGLrg+nxXRPics68dhL
6AgqmZq6GLo+NcZqMqM+/076pTOzLFYodtQFeSSwzmkaozxhm/l9b+Df/4/C0a9U
nFPy09ryH8ne3r68QpE00POOL92QakOkZt76Be3VliFL0tXdkjpEyNSXj38jTk+q
0L9PmvnqVT805VVUfpjfFY8BlnWA6ZlUrYK6dBuRh+oOn6IKbpynjLcOxtIP1jdX
dBk7WT7eJbChXzMK19wWtSKv9y3mCCqIiD9/ewnQOGnggWRaHoO4nxC8SXlBoLPW
UEBs4RGrTTPxxi0GIBXeAZHeKrLtF2Si7yj4BP9W+kHqsmoHPtU+2fqW13Zc0saO
IiNwcCcgH2jZYrw/hVzaEI1yYNqJ5LuWi2yyHw+b7KNVRWxPhECRy3K5tE3gt3Al
aRsN9RKT3AUPIr01USzkvm65zJVYPgdhBXyV5MexzrwKIxJRBajjbnH8C/siUdad
tSBo3LTJNI73uTTnLWYhSdFL0P3QxQCvwv87Ocei0sZMdeI0F5RmzjLPcbeGH83I
RygdsS4DSF8TOvz+zfcmzn6rRUfA1o+s+TuC8AkbjKMQPXlwGJTR+IYVvlW+TN+6
fP1iVM5V8KQtjAUpn9PBiWzzhjuuoNLdyVsdSDxh5cil7Uc9Jna+rURobiRNkwig
fjrvCDfFeRhsH7eS0MiG9ABtr5LDrUE5nx1Nia5E+k5/61yQjNaThhF0/ThJ9KXC
zD+P4ZOTWToZTQqoyLbAdoyspGEQxTgS6W8rMHlVUlOzmlIZ5DJFqciynDYAX4ZQ
`protect END_PROTECTED
