`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XcRygK9L1qHtP1N2tVifiTmVmsUHkHA5O+Lh684K4oBtmy12NuseCDD7/blaa4pf
WsYxo7f6zZnGvsd3FxJQHlYj543k0To+c/EiXWB2lXGcaKW9ltgtVf2VlczhtUcc
BIboBhnFya6hS7p4XeiTztJRHhFS1xSQ++l0qILr/wY7itj7E/1GynVMxP59usDB
nsJDjtxvw+GwDFg3j1TOOvG8KyPv6mNEmGSDE9J3KRUIDfTRpIg32+3TiwyWqYc8
yVggITzmET71AVtBC9hEKLbJeDJjcRF2lDOWfnhwLVCiEl2akpuZQaptjj3NM7oU
Xckn1qWarLylgFJ0BwV5a6x/MzFnR2JZP6SBDycy6085ax+YSJhzX2lORoG7x1e5
3Hqfj3yJ0+Wj9cZDBk2FZSCY9KX/io/DNNEwH6ZAgOS21pjIBFRnCs/v8l0vXtHz
//CXUCtOorsGS/j/678ePfreRxopfxJ/qtil8YfRRmCfxBEdUVADCg/NGUQmCyzj
SW9IjJu7LydFX30TRyVfqqHGxsb1P8VWNLpvO/Nfssm9+S7CKQaz63pHvtWlZ3Xh
CSa3b5AUyH5qfPgDChuP98ZgTo1AIvvARh1rYbrQRgqK/4rn23vVkhltIxux5Qqw
Q/xxnVFRTAQOUB1lTmBLe7UvRWciTt6gm7wPr6QlIF5qI6piKjsMEx9qnWxQ8w3a
1ru7qSmLz2ycRelg0RvMpYcv9Wx6iWSHh6h6g8orjRiNragJL3Psx/ZT+LUzCXu+
G0pOfF+JRiGRH6qIyVBdqmX0R4XcOaSMwL0qbHVt/LKsaMbyxH+kl1fiF7KtLcdV
dfgIOUJvl6+Yvu/3lvYxi9HBfSd/cOuA0qY3ChaSm3zIPcN/e423x4MSY45XQKci
03f2GY20vuwSCyW+XyYKMWjHgUUYimmBcyj44Ji/KY5mcIqOpxQzikX7w1jYbqVi
kslv1rSW6wF+hTEEuAfzd4LKDvG+8hCxW0iRD1YXMuras2A+uwqtJqLToccFzmlh
pHyu5xL0p07SAHUAUDSlePrfN11WBXesq7n0uSzXmSQwhZGCcQn6BNO/gOPN+8tZ
h+Ad2mfCe7wyJi9xhmW09zXGh9WAPSpCeMExDwF64D9mMmOEK1FhO/Eetc3gHck1
GibHW2TgRyonclswJAG2r0i7zrSVGBxp9Rnusi1f6Yqy0WPFpIKctSQktQKD3Ikq
vqYJ3/r6Bv0O9705lwWBRoa9pgEmPtoYN6YzqkABtuWy04zn6jhVAckWR7rnKPYx
`protect END_PROTECTED
