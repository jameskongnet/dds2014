`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nKjG/Bs0c+eg6HJCgZAp1p9G0VtHejZ3YeRR3uTDntyu8vU28veA9c8O+iJDtzUv
L2uhhpUr0k7899DYLkJqTNOsVjZKiYepmWs3lCkaCEpccNTI+5jOCzVRgKi/5DJI
eFIF/3BSWfAbtEI/ukyofNOhKxLd9a8D1n9qRt9YQRsVhRO850yPNp8cdA40lOyS
dNKNZgJtgJLT1+0oWHKblT7Zrn5Vr/AFDEwolkvVB5wKlvI4YZrWd5fRSv4vujo2
fktWUMGU9w15LUCd8jXy5Ylu9eA1hM/ys85DJI7H3lXIiUD+GZASLxKqG8QLmbIu
j4Fwy4MtleJhjseLyOD0MuZig6qIIXStNgJRz/X8sStQWiBmreXxNKFlr25Gd2vu
Y5lZ4RfL1nyYn6/yJli1h4tD92TM8TVkauLb62HEdUjCrYOHY/7RWB1KtKgKgTk/
HKFalovE6dhLvXtb6zaxWk1KqgCd5lcf8ufxqzj850JvUOoCs9d5PWcV/hCeH8U4
YQTEbVm/HsboHNA/lS75SzJNx+33ODPm99he5mRNPjJpriBMG+39/+a2mNoO833L
5KJgU35dlVyyRr16nJXURfDmajQpY9xjVcwWwn22kODrMz/rMcptAEtT7f/4BFUZ
sBjj7nXtCSxJB3/i93it9g==
`protect END_PROTECTED
