`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QvfqeEo1OoD+ku8E84ixSkgFNRvhBGDIO6nbAnCpO8jRTOdvJmq4GR5qvgqW4VPb
82VZPMXL4IzWZEl6ufgs9U9DZ8b9+VeAxQxvK8kc+zdUoESx5bjVohPZXu2OI7Yj
ScN68yru7r57hF99sv/yWY3oancvzXhOZchWiJNgGXmPFt/LIuFJcqPaBBM/x7Dy
3p2kDhiHDeWqD2bbMgv+kZJDqwxorEC5BSB98Rbfg3E7ZoGxw66N5GtVuivxYmJB
5GnnDvt60gtiYxgnvidy0kLnHEexk7bozWWXWvMfSMnoStQg/MU6SsVaeZnl7AdC
sQcK31Lqw/j95TgSk72VqarzA2CKQH6JcSCDEHRe3e6u5JxlyCAcxpVFDUmHbpI/
UlPliJ+OP6eeaZA6oLBjHtSi+LELRFg2yct0M4eJcocsdK+LnTU4rGWfYdivu/Z3
gDK9JxP1GZH0iyodz4cnvH7pGlmToYGvH58XyLCt0H8SOeqljYMGLeGYTUMO7v96
e0dH0EPLXfca4Rjyfz/VqcWMP3WcxAhV/PFI0IMit6Q=
`protect END_PROTECTED
