`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w7LDMHLM7keJ9+j9luAyFpSWu+NoQLXw6OuPn4BJq6fhRYXYH1pET0VErB7iMe4t
bg9OImHbiD/wKJUa2waIGUHkfK35lQXrdU2uuawvMsyTsOZQAQYQh3FxlDx2rUPZ
scdfTivw/TXi9JnvRRoDMerq1XUZCoVXJYRl+DWTLBZF60gfXCozr0+wZo9izYQT
gmaE7qbO5rBjio+cK14t2mhy8rfuz0Nh0M97WQSzKPMta2rmzbCg+gZRvyb9+Hd5
ZQQ/A9V9HKCNZmDy7sDp7LxV/OsQej+QPI1mKtoFGUY/2Lp0AfrXJMO7550guUXN
d6vPIsCacJ1aDH9UU1J3QgFbX2cyl+BT7pIkaF/igN6OaMZUGED3PWTuqxeB7FZd
GPDZ0PrOiEI1aFVvI0tDIXEPRVTQ8JL3/Mr3j4Twh0wkGguyFLru7xDwX6s+Mr7s
BKODiEPVUipPzO0yiiWNxX6OhWL4M826KjS8sfHVANbwFkrsbFfx6sbTRHeVLcUO
qsaF23xz7/QJNieu7TyYXla1ChFva9EqqWgflwmLUSCP7IiEn0HWYfvEZPb2h/R9
WD9XTI79nptiW3Vm4rH/mJf52tjbkqmJ4T4chqaRdRqp745mPpIm4mpa94iOjxjc
fFb5ZE+Uco+PANvSlzjAh2HUzmADa8IYlKgaOMd2eHbaO70743zMyteFQnsyqE1x
TpliNIVNLn6KUfE5zjraYasocLQFUd2QfmMan44yH6JMVgPN6HQ+yHa909/XqagY
NO/xgaReyNycOIwJV4cgNH+kcwdyWOVMKbPngxX8sNH3e4N51cYhHFV8+rE0wfWW
2JmM1KEpRXKEJ9gSEB8r/wRKgJ4GsG5aZ3/z7vbrrNg4OHryVuIEyjN75glllP3Z
vDFX6NLv5NOU8oG8iBtIPeB38jlLDNQBIcdkxyKv80A9YFRqnOFWOxYKMgOm4zkS
u8R+daSqyK/z9rXBaGIE5SjyzdT/LGsxejLFyY7wJ1YP7cCPbT/ekkUeXcJH5y0B
1EkbSi0FPQiCz3EMrmhPDUeslz4Bfasv3AJ1JFH30yv3Pv6u9HrgYLDmUaXZnQAz
5AQ0K2lj9qb3P6tMP7oksCAk4pEJCgqqOvT3IYiAIJHyobvAWeyohAV1wBcrZ4SZ
cG3BIwM9OMFT6Ty1vpeeGxNW/GR49uioR7iKQsi/GzFxHOEvlLyMWDcL1IQHBYdR
la3fCv4Gfkjq4koD9pSHjIXS/hRfzD8i1k6W5cr8w+nnSq1xPz/gEW/qKQUQfyfU
SoY6dyDNTSsNI8PAgH8IlSYgrGz3r1pdZcZeCiB+yAKs9JezdG/FySonjbLy8OqX
bhjfvPkIe+oPlOitchOUdUu9W2hqlZ/PyGFcaB1OQiEZI6a+t6OqennHz1s/SuQM
fYMTbEu60Zwd3MZsyLtx8YJ7V8+oKbDi+tu+MO9KFA0Xsku49+MLFdNuuIBTRDQS
uxbcHIpSr4cWSO/9qCmqdDE+RhIB2kadwckZQvF2Z9a4RTD3da0bcjK3oepcvXe/
NjG8udNexeGe8p+6GxEIteLsDQvOtYv5BSidzMxJPmqhmap5Of5kmCx9BKETjH5Y
PAT08M/6WDhl7GbNAotc9hWDNSbZswHf7PZEd6k1gKGKObg0pXqvG41mKcvNx5Jm
8ohpWsfOditD4HHQpCx3s3wXwDFdPoFoW8481qWG/7KlNldNB062C9fBX8ohqdkr
GAovGKKtezKgaDofr3svrlThN46ClV1XvRrNQ8RLhx1HRr5gsBB5KvAi9+H9F67/
xahjhYY35IVRNoC/UeJ4a9WXca4cQ5OxjvgYOGNA7NDJDX2SNKLF1B/0w+FXliar
xFKi/V60pCbFg6SE8C6dwHUufcuuDD74/UDnaxv9EIuuNZO9vg7z1ISAEq800bDQ
nIiZ40YsHjfVGV1yH06N5KUdqCDzTYyHD2jCriXGyjGmpIx8mzz3hOdoF7YGTP7M
fi3mZ4M4xtEwAu0/xXHuEYeD9yEau4A4MhaG6pwdHv8A/CKdzpJad+c8zPfJGWza
vG+KFlo53VIlYc50EtwunmsfFQvS2CLda6BVDu7mzMu+kRT+otB4i09ckzOKo7k4
CTCi8m9iPjkVI3NFewQ4uZfIDK7G8eOKgDKTSaZH0kqz+tEIy6Ax1vj7E20Uni64
bVk6eZx6PA3q5DzlgegHFRKPDPT2g+g3i4ptDPoy7Yams/RIQkm60+iosE5S+9+p
9yyYhMpiHlyUDo4rkZk+nGqDplPrzxQANGNTafDK03tjsSATxGslRy3QjQQSiIWj
Q0Cjr8JvtYZQhkJIwyF1kSDMfKZQ3lUjQTKiuIItRVeXmT6aBm49pksuRzz9tUg1
3g7xK+KzOrC/8aRPUBT33yVZsjkF8g1gKSwyThMzLZcoewnTZ4w3iJQAF5VO3+oJ
7SEM+kasG2szCpeM8Z39ESDUJyBV7j7ASjodGCIPR4rffOmSCjJGzeEzAhgGFPeu
UfrJC/zu5z5sAu1+mxgvggtwWneN9jijNeCPPn8oCzLZK3A1AmojOs4LkFRS82tB
xSL9XlgkH6VSvsK3qQEnkZNYYPm5qZ17XOjlTKTwKJStcvK2f+Uk2AOzFZ/rnnzB
meynOFBUeXo4ujSBCFyb3VkE/XM/ROHYLzMrqyVodEacrHfHAUT3GK1tEEmiVAy+
Zn51P7csP7BiCyEJBlACMVE8TfG0S1zy7JoSbWe9songnAktJ1gdjbb5f6/xYzMu
nEXd6mvRV4T9M4oKUw2pNBZaSW72NXh6NnMH5qJAqYTiD8UOGlnGwqLmSN2nVDuO
uHPu4gTh0RKQztgVC49i0kPFCLnrMkn6k6jFMmeBRwV3kmELzMC7WSeI+L90s+AH
s3IKm0p2CzlDoVW/j5fywoJRLC86+suk5J6zaLLjImtI7VWQi1zairy00tEaj9hW
LnxFHahXW+INRxB1ObW/I+YAIfZUTLWlKIr/uzqLT2X2pvuwHZ+ruShFnG/iSiKB
lud9q7ZS2z0cid8t1EHx/59M7S0xmhLZldYS1eOh3k/jOdmY7RuJPsG7yB6rErQV
xTcymBpal5VjCmxkqWINIE3Y2fneiHDUYmf5cNDDv5SS7VH0z36b4DHbTD6IGpNk
WaNMp17vsN04g/BvBCt+2JzF5edN63Gj7EdR7AEn2MpGExagucv7fmY68HE01yIa
UDDdqc4zcZFFhB0Q+DY6Num+7W4+XEj0F7sSfA2BZVEDOSuUH8Oh/A0y11Et1sns
ofxuRJoGE2tQbidtqqj8WPw2PFVvVK+CfjOSU0Nh5kXHUKHCUvp6G4ICTQOjYKcZ
5jiP4ecBWQH02xu9ZGxIbc7aGt1vLityTqGO2bK26SHrppQonA/Hqr0SOszrNxUG
axZ4aS3whLexpG7IuDwrgcyBG0++Eq9TaIA29SkuDMe0L9EUzzyboj+Z0A6sd7Po
fNQg7PGCh/332+NIfTknA3nnGaT2w0LgcDA0Xe98z/1CcZjBP1MQArMiB6Ql6i9r
d0YjjGH+1VWnQc/jrvnRizJF4nL5nZCFAcjNZLDsKUjYzLKedfOibbAD2Wsp7u2K
QjYcYY/+7/gJ3YI8nGgMUx9hfaO3hSxVLYlpqy1eEHoRp0gCu3YUXj3xqvM3Epfs
j1N0IklcJfiMeQ4iQQ+G/L+qhfKGc1udOxAiotE01iuvU+bNzoh6nx8xmKkQfRah
iifhQDel/tapz+pszZ/FAEovVyc5DA8EAU+5G8KJZtIMTLcGGO3mm6UmIEmfgu81
RXk/IkyH/epWacw17qmn1P16V1VkICKlfZ/Vp3dExJiGpFcRAmg+V0lbHeyff2Kx
9pnxiBppxd7lkATAVQmoLl/XUt8Va23xyd4Qc2yQjXqOkWK2gB8hh1eMe8SmAL/D
jxLmMNMWuwZsoqicp56FwMioWmZbVz56sB3omCoRCkczR4yJ0b3vp7yQJCUlwlhr
E446pINQQHAjAry7LwHEatiChsCD82VIGC4tbg6Ek0x9gsQV5lFoboFmJQo9xk3j
4FS7cU4xS3zuJe2qcwW9/wbuHr5fb/VjyUKbGwqufTDFK/foX/aLZKQAT27JLpN8
2YRE+eH/BAh2l7GmeEjfBTWYPetKmAE1dtvDVfqLZNHESmd03vJXr01jGF0iBPB3
SoWJf+/Sdu35ez7EQvxS4w61eUqntSY8t3VBSvUIgk0=
`protect END_PROTECTED
