`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRtJpccgWgN+zMiEoGHgObaVb26GbV5pPi09p0KFtcniIarhO/khzWRheFC0BMu9
gbgYL/VbGfcGxJv+8Yw3eNka4l0j4GVgkdCzAWmoHsOH1lAzd9r1pBeSJWljBwK1
hW77Sw6Ph/WoSW0LsJ0Res/WD/9YFrBdegoQ/wVPgyuxNRREIVU2OMEuVP1Ue7+e
aLbQMJt2xrU48fMV2AF7BdfctIi2Z6gCjXzNsh0Cfb8MDRMUJ67iURKfM+UKXwy2
kkpo6CAiAHot2ukENe/Rc3Uc+bbYNgX5hwXcVVIWoexTWLOBUdVsarDbFtamTYuF
UbysFMoHkDnUEZ/FKhPsJNfvHhVWIP8SIZHDvklFIfxBBraVxHq5qfXPagDnVvb0
pO2QmIobBsYTJEMUraEKGhDG/r1tgD3EVOFKenO25Lnu6+p5WM+b12Wp6VGADweF
KSeqJ18d1MLoF23/Dtx7Nyf6R5Asg3+IttoGLtEDFC9bKJGckl02tlmozoFdsILJ
0XFpxt14ab9KLWSH+eL2L8CerE89eA/oAqJgGIqMu1Hso0eAgvRaRRopf6bgTYAq
/ttbPMCsCurtmqZoaMdhakHz/HxyRDTcF9kuJIAqQV/33GRwdixz8rwsubDhHFEV
jYwAESKPnJ+FF46bP9Npa+ap2VWvIdIkDqMJlHI9rLp2umnqT6TlzlJZv0durnVq
9hIJL5nWckw8jur/KOKy0QSNiLiQOnq1PneWjBDD1TU=
`protect END_PROTECTED
