`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I0R/fC8EnMPV2btjHUUscI7tj/EYNGv7LeLRw6lgEKQoiD1+xCWPA+5MQ831feMR
x91yuOhegd4bwIg1iVHkKX6eg+EkXe447ev73/rE8Yi+Ib2LEJ3ndyHlXMMbdJKW
PeSPqI2SrndIsuQaAl2u3Xl/9LRXItly02afjZWxJcX+wLXAK2dZA83LvpRH5wh6
G297eO3PT+AI8rHHXRxfvqI8Ol2Pq4h2LXvXUuTaXhlelx5NNvjjoJGX3xdDP6Ca
1Y/6Spxt2JUwZ6VOgX+NmAHhiT/rqF4z46UDehYsbd8I5TEjFf1wP800DSdISt7T
kpPQv0DpBkV9hWtnT44KayQqZESCvW1Euhb7j6wVerRa/mMEbSFanpMTObq9MG6K
6yCZ6Qi1lNpc7RcHGy/Q3icwESZMyoyU6xqHaf8ji5iLXC7Eo3h+xZrEn6iBROV4
SzDgJjrgCsuFxsxByOf5zu5/G3SpB2EPGq2ISnocXk+KikFoFHbY0qibpWfsSjA7
BNQHsk+eCVjyAGWHB+Ij8ODzAN0hWaX7k76f4F/egO2ZquWIddMoUpPoPD6uoiZ0
GuQFDq1t4xhO/EPKECN5FVQf+b9Q170lH1+Qn8H98ab1L/EEYlO0i5itYr8+fy9N
JlyKdBGBwMJgqgLOtJeBlZIQXd26sS7X93rZq7W0fAD+LieaWxJWps8Pk/UP7urT
1morbu5oq1J2ywDTKzoya5Bzqhgw5UIK1AqwD3E69y+2DLDfkdXwURdIfO0JIVRT
/jabHfxSwoxam13rB3bGhp6n+ytzN14kW6U92I8yhkMPCPM0KjD4aHdN9V7O48oQ
Wl63ig9oFH2zufMNTTp180p/4xklyYtLCJ++HLsxRnzdgbKv8C0EYLv3VLNkDy3N
IXg6ofsYrB4sRYQ5smJmKBrw19MqGtupYH1cadbp2ylr0xb3TDiK5qxBxE5EhQdi
Rr0MjAZmQkb3qav9hFsijRU41CaUJzDZGzNylBIATBJ8Cl+DYdG/BN7ApJHaSMdZ
vyFSJElUIlVHELtlfF1D5tan4f8cKViUwahdV725nETXetMSUANURXah5/bb5eh4
RR7jBDNASI21aUsPFl0XNlHezawtF8R7X3tQ+8VLJQcX2MbFd0hoSNGDeOQra+s9
QZY/YD1aecEOuGu9t2asa6dJfVp3lOR/ZNFXADwMFHifl/81No1FQS0gXY7+RcrS
jHwcKc0wFI2me6U7Woot6bjxpV9qM7mLDywmd0DtKsZrc6OGjDv5ZfNEn2byRXcR
Z3xuK8WyznOWy0Hdp/g3tXdOeJDw/g2Lzmww1FjHUpswvfYksm6JN08mK3ENj3ic
piLAh/8ZAOn0jUDY9h9Cht7DTxkPh+8/mp9C1TdD+Pv1Xd/TEnWhz+vG6HGIM1uW
HbnKwo/ALEBwUWHQhMNl35nstMWj0OUUBQR4c3vhCkiv1X3uKD0uVX80WSsY/OFN
7RUVx6FtEGjYaygmzomxxelNjqs3FiQGu6cATjgAGXs9XQKTchAgEjRz8g6KRwur
cLW4F+jPYVxnUqFsbnojJwO/D0QD7tQUgrYLpvb+MuL34IU2Oj0/QHS6d/abnhmv
13b6u5Dm3KIVDUygB2UJKlY/TQ/c1aT6QofzSMPlJdlaeSRAQavb1/4Ohw1H0oSa
pZSwZsGqwLGlAwvyNKXhUL1Hun6JXgdcdCk08tIcHGAa3BT8rz1HuRSjHDtU0rNN
i60z/62x8iFfRelLn5vVPBRvmE28DzRfm7kZga3yNVLAjamUp4kGYHbRBERS1Hof
KBCvu9v0JKNVeH9QIz/41Dvr5AAQHRSGCcCsnN37yiH85xYyBbvQPMXObvBjfNkE
uJ3PSEbjrTABx+TF6vMdDJZ2zmDyl5KvXS/esOcpp3+li+Zp6m08DavteQTKV6Bs
u6h4ZD2Scl8eIS7Jb8CMkEKdOf0EeDCjYYbEzfw2lIdEf30wmTiWnS/frYZqcF01
1Jxjq1gTqMadg39BYI40QtH2n5XW1rZdfG1ohgAjBj7UtpB/Ms2Z7TTvJvRcbWbC
UfHyxyMPAH74h6a8/CuxFhH6p3xg7fofpTOSGC01NZb7HwR6I2tBKnTfb1o6/1HU
XG7G00cyB3njpyyS+owdS1NEiqHZyV3GvSojazWrurlr9DySI1ExXg6z0tEUE3Nb
UiX89DT/2Yp99Ajercr1vASGrKw/4qq//bO4DjDMHLTB6lseCsSeQAt5lKfRXTes
x9f23tTj12zScj8N/iHIeh3fBjjAABS8/7KF0vAxSJIa3/MB4Q34n0Zp8P2NXOC/
Eaz5VW6ZgEgthwjV6UMrH1ARsTzBYFGCIZe6nfWjqeB0CZrJkTu4Gj8k2GqbZKA9
Cg5YMdmB/98oESZjA1pSiD7pxQOMomlf/7i4odUAN3RhhrGIttZ1XQPS17jf0rzZ
PyoEKMmTAqQAJ+KCHZO+MrWrYp5GuNLRdbSJEVUXMSRGDIQebXNEytNrr976sUO4
1zwbupUCQMU4NftGW45MRxO2CHnAb2NxAkQHP+Mm1cu+mhg403/Iz3OE2eHX0yQ4
Ub/FQ3IEC63WpqN4JcT7SX+Iu2QGUANnfw+gdPb4Yym9FE3fu6DX5WDFpLndgK4y
awYfrogvpmPGKRsvFW+Gy4fCkGyFWLXVr1Tg68aGbSvJMNDNwOxIng4Sh8qN0HkZ
S1JoIN2sR1UTq6szcTh+C7gHwlrNfrR4ue5dssyIPA+5lCRiICuOjM4Pt4lgzaQ2
IboudTYc9WdvEniGRbR5kkvl6q5txE/ZRIqkL5s2/7pHhmZoxkBuDjnHKmUnHkHh
PJNfCqoiwAGie8v7CEd1b2OaWVshWEMBUkmNxBUms0o1uBvOSIdfC6wuPNq01/yy
cVGB4JNkUtaUaccHGDVaaU31f7pgkq/Br3vVBCP0l0vd5wW1Z9+UKr0kZ6F13GUL
bjuQoLi35v704YSboe5b5NTcJ0d0/8fjen/+M87VCS5ZsAMgqua8oICimpXPN6CF
JxrLV42VZu8GfmFBNoStMCpUNB8/Jd6EJh8AI0r5sWKgoTRXC4VNKxnVIZ8YknuA
ckPptbsA26X3t3TNCWJRtB8RLF3O1Gmxu4a+9nkcBLOTXeMc5rsuT4V9ZFHsL9YG
2xkgPjJWtu/KEizO6LTW9GcMspH1PdJ9aQ5QBbLXSxYR3xsU9QUfZmtJMaXlN7lo
TgMfLu5sTz4LMAGBzL0nj1YhVHIBRyohaxXOq10N30yvWRirWDG9rhNS6RqUVruu
JM+bSA5Ro7Kv+gZBjrVStd+GSx+0gFpNs3XzNlk2XZYhiBRSwCFsn33+E2MlFc43
OALgcp+3rO+LVFYYpcrTknd+ENKmL9tM1GJXkuVwy+r+hzMTNys8YJqxYhZU9oY8
Px/eOGC9zIOTrghx6S9LFGVFt+vzG3FZE7DkIvPJ7OLqoNwYdTzo2RNX0D/NC1Ow
vYXnQNJLn3Gh2iC3+peieZUgZ8e/E6uOWIiaD4JVb2xhwYHVbCaO6RSJ/hvx+YQX
/9AX4XYyERzxKfRrh8F3kZGo2YXiOuqhirHuFaQ8CzFd8x+i66/dV87NIUjy4Oxe
ivflVxMD8ArjpIoIWb7rsTVR3eICzzEYbTkuecU3wDtLrYU3/A1jH6sRjU0TXDSW
IjmDdCKK308RvmjdrtT84LUS0ux69ROZguAwxed1TAWmdvdKEw1+Tla3f0VbHDkw
SSgrTV/uHOyl00OWw1IvLQifjKL9nZxZ8sTfIJlRn6KunVVN2IXQX9PMY+lVxKeF
ZsqGIhjbdiQOJ5itsUbHlEJJPWJmw572uN7E/7qNQW5ynMF32prjzs4TGTDx2oMG
QUoEyKfh7eELaOr6euJGSq9S7SB41SrbFqpQ6G6+/uwFLSdTE84/n0LJhLuENLhT
dIHX/t6IpSBkuTJyx7of7fsQuWZuci9WuV80xvTI1f/8LI78yzb+z7dC+1pqUjrQ
4MAlSINV/IYvU1OSTes0NZpAJmqHyIPBd5GEtgBUL9S0YsvO4yrqTUzrHM0KRbm1
ioMdFRFYVm7xUiTax9IJae55uC2YUYwXzgSmc+FZ5TX6LPippbEWBMfS2p0HoHUy
t1xdVC8i9H9Sdek0DYK+wIhzbO+iqbho/ktrdq9cCM5wfMmBTrMcTfwZ15FmRDVj
dTwjYTCCWhkVUdnr6uEsy1cEMmJpTbvT21BR7CV9yCu3YQqZ0SgCkiD0vZVoxA+L
VW21A5gu04etVOlDC3u6LmNzV8WkA1+A0YlEFlNu0UowXGQwg+xjvZoal/nLT/JM
Haf0tYptgBAkYdW6j7cXQe9g8hIVXLh1A4j+tD12RTaoKXgyeE7U8LgESuVGJLqE
BSOLAddJgqkbPZDogofMIBeSPm6MxW6Eo5OnyKDv2NCQAoMA0EXB9YkPHCwirv88
g/qHg7oS5R3ZGPJiMPtEGm9o8gh0BhPf2JzlyYNOF9zBi1wqc55ltCFsMe6NKD/Q
Krqy/sC4ZbDoxk8UoUNeTGuCZqdv6joPpFu9dWeFTlXMgfoxzYZceV9zZpGTuvmV
5CnfNXExngxfezWu7Oj1toboz0QvVyH+aRTS8PBiruJAvvdQW1jbJAQOnwVzNTFg
9woEKH2GSuxwljp1porfNKlXKEr1XjoV3D55nr9kCvHne/e4m6Sq5nlMoXdEDwng
2YO7/9FPeqpm6DGx7ocwper5vIdJlQqhG2DKiD8ReQmPXGE/FABnOHu7U0RgCe/x
Z55JnCHF9jM/VHJ4YvizJyopfljMZYwNG1nnqGoeYefvo7Q+Q2J2pxL7kmVqJjNW
4cCgQq9yexWhmFwDAhf8eC/OnFUTGmLuBSMcpu5OxWkAIwBXHBqwSTwJRRY/zpSf
RnseaCVcFaQWUl/Vx+jkBlKQpK1E/3AVHnfB8K0viLpwE1I/T2KCDbd6851Fx1pw
d8ImSA+GDjm9dVZHqWdA0Srbuo1sjfR4r5e8CqWjgw3XoVDrCdKoYmxrDNhkrxb+
75o0WQj3YhWXzj53TzhgDVs6ok0qPVVkIOl2LaXdutaLpPEJm/K7yRHlYS2IK3xc
Md/x1dFmpglV6lMK9YOO332YNYuF414GBDzzK6I8QUGPVL3qqxasCelTmxfQQgJ5
rog9Amh4lEp5uqt3ZWXlklhK+7+gH7F10vURtmEs98aUXN2wdGuF52IAtGSxD2Vx
L6/3ouIoGxCPrTLXYXkMmvycvOXm0lGXeyjCFttQKmFiymk6nGhaX17Kqd4lGyGR
98p/rGRsoNw5AufhWeNSV+g/hzGoOsP2ZjxdYr8+Fy7zCHs9/jIQkAZ8+RoZ6hC5
W0njLFQoCrhKirngsw6JH0CQQPy0H34MJveZEIhLe8L1zy5EOscV6pYmTWlFRTdv
orAnac/PB40FAMo4Yly75AMBMWo8N1geU3l/pU5pB3K8jwHtZiYls3IR4te8V9jv
I7DSAM8sj8EARJZIEUy/aYLia2MtnYInkY+MBhQXzVm9VXJ3svkNjnVZTlULLWQR
rF9dqMVElIdgQa2uWYLigIBp+aU3MqjZnzmCNjVDT6Zem7fe+iFkGoowkrt0Pxlo
7JYGMMlaJbmS1m7PteTOnbBvafzwpkJPVWDYAkSJ974gNBzt2450DEF0TVa6Eqpj
4e4/s/pNE9xtyaEgENgZRb2RqM0hXDdeUS8yToDXTcuhRxw/1oKZ7NfbM2DZsjOK
2NAtd0+bri1JYzOx2v8kkpMfvQC8/V3bytGQK46oFQy4h/FYr13GNGDbc+DcbEx9
uTKVxZ5+nECClB7xVruB7ARJCyysCibXgY2A5d8HiyEXzKYPmP4YsSQlEsGGa3BJ
R9kLvbvidUJ0tM0NeIDVmREG4iRx9PyY2SPxl7/3Hu2s8l5gkP7iJMeJeIzhfNdW
8R2Tdx+W5nWMlS5f0fPbC3/m80ApdY/6D8Of9m5Jqhy/OVoFI/RPWbyKBbm7q5HJ
FembKeK7n9/d5a0v5ivyTqsgnd+RxXyLlcxjYGroZjFcGEyqqjrrJmcnCObokzRz
VlEYcHnMCtDnCBvckO6f10N/wM2vQoW6HULKs+WyO4b9mSyz5kRqfcwxDPUlUtBl
29Zzh+JVYdT3xYURE3Dy+vLSc3P9mOdjJtU3M7o5STiJ7s4H5LxY5MY2w0LpUdOh
i4ATMu1nEEXW1IZEw0/3YzmwumhZWb0ZQeA+6mT7ZF/iueIdbWOFTMGIZTT2AzWF
R9sFC58eZyOsBxbnbt2oYI0NHk6DhSJk/UsibQO0A6t2zO6wisCeXNUCw9hOmKP3
ztsZ+cVocdRKHlBjMgILw4cdGYdJJhoDlbAyChlK/2kedM8PbmddOOMQjbFo0nlA
CkJW33DAPMx5frGBO4gMRwyFjajiEt77P+521bJaDKh9UadGlvD+O6varB0uteFr
AAahmG8rsssiuZrRRiHDpg==
`protect END_PROTECTED
