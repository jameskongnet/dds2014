`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d534TlZlWNxfboDsZCWZBSb14GYD8P7dL4yMYHr66KYgGhx9QozFq2rX/es3IflC
dQhEw1sETNywlHGaE/2NQmJDZIcPM5hmJf/DWb15ajcPS5SDbGEI9R/O4wcAtucf
cemclP/77/9LrlR23/ZpBhELTHl6q64x4otIp95UhjJ58gFBVTHXnyTx7F/fv4/9
qx5vmZnXRwHyhcXwxkUPgWhMFQZIBpsYaqfaAS/ozDaeTxbzftIrnjOS/1deEMc5
X9Pj8QCmsekO3+WrCr58qiJfka03tQ8oMm4uroyFMdDUrcTm3esW4VSihfmAyrcy
m4LPiBVnZ1twBrwIu6Hfg8qSC7GG1KHiYQOfvXYOiw5fDae/4kruO1BCg4NQLrSR
l54ODkyVxxwE0B1GflBTLN4KIKI3pitR360WuewmelATFnONSP64n2x9/jl5y5Hu
4gxkkTJpI9mhPaRe0SlkUeYMEZ2EUX0JNWSxkbhaDLl0vXZYnZ1dDeL/p4DkgFiE
v7k/n1erv5Bjlv+N3Gi81q1MQXA/jak2rMZmHvtFdkNa4wfM1ReUP356GD+pmrcn
uX1lYF9ezAZHLPlY2pzlUflD9roob7jFte+LpISEQr1QDMM5R5dWmAyYmb2ZnR6g
0pn4BBQNSL01gOT/G5Uag/DrZjOHFE1EbDHvFtJdrAURsQTdzFBdTSNdC0VEKBQz
r8QPufBJgFYvAERHnId+CwEG6G2T8RFLIhguL2IcmHEbBW5/LIWdOQePRd0mFTBQ
hLJ9DX/FmwrAxjmDNcxMv9wNwl1t2QEWvhPvuPIKMa+LwOHUwcQU9DG2GMYlYkZ/
8lsRIPIRO7IbIC/ZMjn1xA==
`protect END_PROTECTED
