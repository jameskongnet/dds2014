`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wrpPm4JxyOw0sxDocjhlEJiYb8lgZjpuWQMuViE4z27AVVe4hvtMYvJDYe3ucmVs
XkJO6helhc49SwxVGY5zna7PeXQBNXqwTE2vqJbxb3ynd1PsQQEE57B0TnpyCW58
Hi++D1aU2t/Zt5UPZX3A4hA3QQDbHlpoY5PylH7RZVjvKThb9VpBBv3VI2hdpGjW
p+IIgPTdrlC1yCc7j8iyjNdl0Fsg/6cbaW/qR7kFuvfzFqyj1vStSyl1KUMkEsAE
IOG8KuETMfoir0hSqurWzpYhyzEq/d1Yu837OfrxkuDTHLNJ1I/62YrfqbpyRcMO
tZ/eMM3XOK+rvIjXcTZ8fgqrTgxXuwMomSWznJnl3nJc6kMejD87+IEwoDBjQ7jR
0V1rvl9HYXsvcX9IjpgG880O015dSt59f25JksVV0ylj4zod/qDU6xVf9TsmSCtG
dTo4wFzNByt44wIRefm/bfvx4JXfpUy63y1wTdX3p3WGBkqDTqhbWfsz5XmIUr3U
IFI3F+gBc2RWR8sGYCxdHCgui3MrVvcaQZiH0g93aJoc5AXxAS1X02mjul3LbMOo
9aSJkq2U42zzVwXXIOflI0juvZHZ27zs193snWHHrTMYaC/pnP6NLRTHTcGkQcrQ
/EgYfbORVtR11Txx4oL7HFiROaMcqfZiD3HTcWOi9wUqw4TdAeHh1GNpcUnHWElp
0w82CGVvzwtv6nXxQzKmMXH+ewbCcOBqyDVNbZretWV1knNAljorD5LSx8G0CkwC
uDRf6i0YnSw5CP49JfGH6xua3U8c44EUpF96gCRsEr3q2hIFmqC6iTlLs5QPKzm4
eebiXLmeiM/CU1YpimIVxw44IG3Yf3QSMIgh/qGuAaBPQifg67804zrk3Huq/jRm
sGqMnbJLNZwtLsKh+NBUWth0etwxtS1pW67HAqaSiKDN5Fg4XNE8ugpkU5QYiAL4
lBzwDGVfsoCVRquE3F2oH9S9qu+g+C5nQewpd9dlqNP4IeOak/Vk92Qj07a6KMOg
bLSwifIxyyw8Lw+FYbKhVuXhdeAjwa0/AINqAiPmzZFtEfG7eIrsSZ8q6aNxfrLP
MHOVdiY9jJJGgSYjuHmuWdpd/oLmfKHPU3RK3XKMIZyycXaAuxGIJ+u98hgWXEdw
VUhnbHAON0bO12lVF1WCDsqR8OpT2HFdRsDTpjF6B6ow6BmNuIQu2Z2FjkA5m44u
Hk0Go8qbFIdkVfYl4vH1Ccp0unbCgs7gjpKysivk17QcDhllcOvWtvcUxGVXjk0K
9ZMBfxGaaYwGJaWuaUJ1kLhgxOIEa1E6BNhR9Z1yr+Vk73y3fLoTG8xVlmxgaczu
EvQY/nAoXZ5L3zboxRlbUOkk+59cHjXqim4EdVXqKFIRornYHbXtiGB3iT04BZKx
QqCSd+Ju8CbzQJScj35jn0naTt9wTe0zH/yMmYycKnfgpLagGmy+LOJ1QzLyVFhy
cSQx4I1mJJ1Too/6KebvGKvThWLl85sQIgjMzds99yYuqW/4i1Yu7q/zxZKdiZp5
AhysrhHLYhaE5dpMJc1msMsQjbZlBnBHyogOwOlvQcZDQsFvdgGER4eBo525CSBr
m++i4ON0oMKaK0iasssn4BKbQb156zVSGAzhSzTobIio7EzFAgJ4JnO0MfRH3Bgh
6jXukyReD3ovfsmmIMi5W2MWGiRIJnTJV27N8lDIUVfndnPWnFf4M9qQ+CFfyM9q
pOWYvx+w67FfhgnHd0lJVUkoVwHp2x/NYN5TYTPUTpda/7g9TiCvVBds82BXntrA
468Iw63IGEIcIovNUNpRgM8nu88FoaVdZ5ngBZDFvh+ivBlf9Y9Nos66xzkCLqam
1/4GCYajqYCx/0sYro9rtIZquSUQrP9U9kvOrX+zyaXMD21cHEhZgRdjf12UbKHI
oqYhlYfOboybVAUYfLcgbea9fdg96xjSrAxtfTq3chz+bOZMk6Y/LTobwXy3IMHL
nBSw/iY5rL834FOFOzbGn/UOKh3ZYTN82DV0lhGhUJ2tlgX1RDcBlOwQKU/ZAySP
/XwjUXQM+4jUMGCwz7SqJ7UlTqQRHQwQrwPKGG6eKhbH/aL6+uSQ/oExi4hKoCux
BK9jNrIj6QBiIDVqBSicKLZsVUrN5EHKd7bfilobi4h3DICgjBRKAfIDUCMQwYno
y5bnqqyE0EHDuL6LmjUpCoqxY3bne/MdLyJ0Lm+iuE40qHuQMCn1W7+IWYy9OVoN
MsEZNvMtP/UoJuiElGWWX3pmWmc67m/7i2ToJrOEwPWEPaZDk4w2rjd/yfZWYU97
gJpdulYMXyGLxYoMpNZqpXC0Nl8IE/kBjoXKmsgduoA+cFIGD27KXJNZb/A6fLxB
uiRBDIoruGy/nWZgZvodCWxfWWwPQyLFAxzrNvsQ8hZvT5SUeB8OmDaRIGzeg0kI
IM0JZJhVA9fruAzJolbwF6B2MnDswEWdwAXD82jC9HqcwsirphQlhzPE8kqoeh2u
jAQsbh6qAs7CfebPkcpyVZsqAcyMxsF1b1ZDTHPvRy5qKwdIg4PdQY7d0cY3MSOM
zIbCIceRBTd0PPSrPTpjeAH+Jj0PswcBKgKubtj713H8Xqjo6i2gQgbLbaJvGc0K
D5LlroRlHVJTCSbBT5F4Z3782IRIJa/ZMy0k+swlVdk=
`protect END_PROTECTED
