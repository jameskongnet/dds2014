`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8aieNjWEx3EoyzbJq49/38OfVZaOonFDnrBTncczoUASPC88vMHky9AF+2/X0+02
KPKt/wa3yTpDDp91YE3Vre/I6IhprBm95uusiJmD5QFpuUkOMX5Ypck7Qb83vYaJ
H7qaNtD+U9O41B5NJ9ktlg44pUBVMbWAMdOJ2sDTl6PB92Fjv8ZA8ggS2fxPLV93
sEde6c10e3BTejI0o8nGJIZSUVJgJMOj1Z47IDqsGitYkITAmIK0OweagVsx7TKR
TIIVYLl9oXbpP+l2Xgb10m0y6H++5pFl83/u2KMH/rFb5YTYdynzrVzk8EnuGjag
kWLzLpwkuxFsRMeNeX6cFOF9iOpxMrCVGY9kUR4dir0e9EPND/EFwGD2VUIdDJgv
eBdc4RYM3LmK7idgE0NKdIn+xOKQsFVjR9JbtJINX4TxgRv9sOsL9fv4LbBbz1x2
NBCdFrOxHddxofo6SiPMGoKrFTRHgn6vvALv+6NJCBwc+q8slgGzlhAQ9sWPc8f2
/kt400l6gamRjxKJ4NzNMa754f27bT6zY8updMzcqi0Gg09vyInu3z/auLJrZVva
H5HwBW6UtQ+BTfZU8VHKEHFWPSf2XKH938pZ6UO5xakW9Sm7ZQ0nWQpvfxCZ1zoL
WlJ5sOjsV4nP+Nf2xSwJx4UIwCv5j7yKDHm/3av/Ndwz202cWliVt+uuOkQGJsS9
77f4xWWfuK/EkRCuj5h97Mkpu+moX23M+G/ptsH8y8pcV7wixTjJY45620FsTy4c
m4whzrvI2A4RonkCd9Mz+OGYsYaDXLrq1FvU4yU2wLNXIX9XWuUngm7QWzAyhn+s
`protect END_PROTECTED
