`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VbTlA3ZINbcD0rdAn78Y775xLk34ydpsEnFqeyGHNLufeq6wjVCy2Bv3uqvQv30j
wDCwfTa0PIi307ayIRRDDMYGdGplJRPGh3vytNYNim8CldI2LKDVmjWgPCMG/zLn
JsXtQBIFUKdT8T4+ZH5L7r0LE10d3vNXgsCbNclewepV1QpAa+Qy/dV8rmxiY5ce
OYU7d/l2UsEQkrHNS0INnglkYaVjMAJByO2VX2yPXuGnJJlcyNb8F88tFLOpzf0z
3XF4mEMG9pfnsXkA03sMf0sNnrOS32EjyZaBvyXxBfdhU1ZtFwiaYV//2uIwgQvh
yzGEFnwZC4/ny3dg3S2q7TNlEYkaarBfgnjKZ3kdb6mvHJfiiu/Fs64W/o9KU45t
O2vTEU3By6B+dMfWR8fpgf/mLpHSGzoPr6Y+KvbvJwmEW2SNdlk/zaPfFVPzfCUs
vhvRlYsb0L63IH9bCjm6VHRM6rA05uVDMDxTQWP+vvELFjLtN7z/BwzLqJMM/Mdt
wmX4wSqf00bZ0lKeiCwFD5DFwXzlIQbBVo9uTtgsrcRle6c6NOICW9+Xp0f4IxXw
v41fBr5PjImprUARn9c0NWiJCsEGPwt+RNV1a+RMI5Jhm7Rj1MpLu0CGtKNfZi08
VwqAa6KSWlP85H2ymLsGzrT5SsZbuX4GNRo/qAfDSoBbe9p9iijDkX06TpJeM8LA
VjUTUKROCXLLxzsb145UFthP+/G3uf2aUH2XnRiEP2oenL2IKRdJHqFf5JEtW/mU
QI98hyZ8f2cSk43C/HqyXuMc1bcHR5ZitOgMbj4ctDs1yq+U29C8ODcNuQBpxcSR
jIwIgu5PYh2p2lKCKEdrf+bnaBHty1VmxTm0l/KtHOoZZ0DE9wziZhSh5fu9COWn
ErsTWc8SB9+Oxe4nw4r+/yWWg8plKs97j41gzgDdWTxOsBG2/npA6mM0XK+rlt+/
bbCkRwEDas6xHxiq9uMrdWTx/w3hh4asC+GLRNNT7rzYfcpRJkdkieBken5Wvv2N
mEd00n7z0Ye9ZbukGdVEQASSzDcfMSNY67d46bn15LWfi+2WiQaNNVVM77AS7U4Y
ToD8pWkHgclODzIb18QehsYfY8imd3RSmI1R6A8BVfxGO4rDsB5FZ9YDqG8+1UwJ
C1eS5vSxmptPtSqhCXcaYda+zOxYixKEzx/jA1/oMbws/8YrGC2NZQXzoBdovlLW
y/vWowiKJMr05NP4mgHqA4PgyK9JcohivN7D/emf6NJrQhPWfq9NpV890NxKAZkZ
JZs53yNsuj+JQpRieGHaTyEEmyz+7zy8+3BuzEvNReh2P6UdcRQ/pQoMc1s8N3zi
O6zr/RXPoYQQ6IOBQ3n99c3ZDCSScG+rWPO9BnDlfGAoGWEEtFUXZVnRoRL3ginr
Xi6pRrhOMR4bHMUlMohPLvsiU5EOS0V1Q2YBzizsDhHCJVnO+vLyFgjUK/OHVbn0
FId5xRbJZPE8Xnfk0YXC4r0eQ002lxuysvcfsrNXCDzS2cjrKL56vuGowwlzGVSj
LO9DsdW2myktVKFu9GFRmUzGhnIuJ9ro77vtDhqqQnankN/EzX/RUnOJ9i9b2jrT
VRHPiFgxXL+DSz0OHeIMAGLnkodGwcmd+45AhBiwCs3yDMbRdxrlEyr/vlDURjl9
XrkAnriRP2OHrfrQHLfooU7k0LV2lVu0WMEqYNTm2TeJncOHsbbz2E2dvVbp8AuD
/x0Qm21RxPTbCAHQXHUXc3kji3QlbjZmHWHPYYrEnLCGXScurs43/N0cR/oe3kWE
BU3qb16sz2QcQbgKHhzNAcVc2q/Lyn0lJe8JG6TGbxk=
`protect END_PROTECTED
