`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rP76GQq8R38YzmRV2cvfmsKbFocfgcPE6BWWe1lykruk64jXBX7KQutcVV7cCEE5
kfeWuKX/g6NqjN21h2+xHZSykF9yWG8RE6lXGaP6kYEhJWBENtuufu4xLMTNmtuD
vJL9QlPwg6TqOlasFqq8mvFt/+ehaR8L0Cy93NbYmZtOSHsEXlLukvp0mHaQh+7j
H7+Gd2NA/ok1ZOyO8FmNeRLDIVNL/p5v4hT5YNBSRFUXD/SyL4rI7w/2Y+kxi182
FavsRTU3/FkPdUTr5kY2nm0iD65opPAP2c1zFM4/YxttxtOdwZbNYo/omVn3r45T
0w1qHe1hgeBZPRo4T15cSgVHvcJzkm41rrE3pZ7jLSykcUa9FMjMJGVNeufx61VA
w47difz+wvP3IPs72Ww+QKoA0QzH5sOC8+uA9n7TjpaSHb8pBtqL/cB6+R1Vcu28
a3k3rR8+HFpTLGVo32TuOiBFmFH72qdFB5MywJCgJoQFFilg8dyZL6/W06F3XxSm
ON54VD0h2NXbBNv0fywaqwI/7MuQQmsJuZq/Wp30AJh8wW//LSPfyrMUkPFLMRyH
4aUTNxTyngFZL/i0vd/UBOXp30BvbQqEXz8Wmv/NPSF90UpjSM5iuzrIemHQza4j
3Qz3/TNQiH3hMHf/RsqV3ixs4QnRl7XmFU55DUACE4ZQFdwj5+PA1ldU+NzUzUIG
4gmMPg7zrrhu0PvBm18OThjxMOFq2VtJVzIn9DtoAKPdtdYGXZZCon5SlyoYpBUZ
fBvvkD3XZuzwos3rXTP4dTHBnAfRni4oSxQj0sdyNqdvNcyBBqZ3NaYWCy7ZBi/H
ie+ypCtPmHHt8TWHCKZrG+4PARJH+3DZY/l4tn3W4ZM=
`protect END_PROTECTED
