`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oD5V2iZycIczQML7kflRA0BdLKwOgiywNXSNu6VXr0PrG9KHc0J4GMWZkwjwWCAC
NBkArZs20n/ZbMtUlQqABt+WaIq/N1zIYupP+at2klMtNPi9UMaGGnpPHvLOODLW
jAxkmk02QIu4776s2dTPHYkqjo5p90tjIsBZRUufNUq6q1MEvPvle+qkpy3KUerP
Weq2CSpWa3Y1NE96OdhME3RZD6kxgQ1lN8fF732SytG0FA0bvuc8aLmlVe8ydyC2
IdPr1rH/UmtIL+afQDZQlGTpw5DJT59gAivSaAbqdQkUNrrY6exzV41RYzMkTcft
xOzSPCk4WHcMUFu69Nx6z5sN0givRZnKdorK1KTWRLMRdijiq5frcSXU8i0Jz9cQ
y9PPvs2ROH5A1HtHsD7qRBPKTNXwS7zF84H8goxP70v6XR6aoEtVwMn8BrZAuGLE
TG6VCozX9Yzn0oKmtXADGyIXLnscRXF/WafAxU7rN/QpKiHYwGseC2ZoTEEDIpFp
Lmm0Rz4bteR633NJGMKnxnHpLqbp8VKpeZxoleBHOj9kXXOlSERimmoED+0kczBY
yYtIB2J/sFpbFje0U2jTnPnLzeVKQqd5jbUArJk1ij116j7BFQcJjDVkouLNjRCP
GMFJ34LktVDV8TQYtNXzbrD2vLt06nNtW+yTpdy/3DWzfQo4WNHwX0GwWIfjGE7W
espfcSW/GlgffiZ250TvegD7u++sQljXZTPGlYfUajCejrtilffrjJRQ1kXe2Zmz
NgC6fEKHL/YkVacTmQektXZsK8RSh70gvVeCwCHh163Zf0LfzP12n4RpOwWSMmbm
K3fSQ67EJkJN6Wgj024bErGIoGkk81rRbHjjFgCu2lYlhzSKXElC3KR69N8GO7Bu
gBbrF3IhwppnmUS61IXrasoRLuahKm4G6nD2ZzZXV2DsPDvJzgCgfyxObqhbDXpk
5ygvJ2UX/QzdUL6HbHKB1AVCdsaZKLvNGbXJ8+YTOxdktX2YIY5QTWhxwxOzx6ON
FB9FTfbNFcB8ydBn7EZ/KeEoLdSUmwP8hBbzthIzOscXgWblXOyd0GZhEDl2R/aL
lCwm6+I40rd6PVIcZo6Qi1+F8u+XVeUVEGJ5K8XoaDr6TxghOhqdP1XM9i5Gx/lQ
n71ASdNaTjHRPis1FhaCBgWOIeR99oSk66PtEEceN88wLZhKxkebveFBJdJHKviF
aHvDSwJynlhHzqt2TxHz7vL8M9jx4dF3oE1rtrQFsprBHPxy97nSpfrg2Ymq5pvu
quknUXmLjpRKOVlttWAxkA8t63IDzXiYB1sEKLNVvyA3sYNw81j1kUtOOqot6JCb
1KCewEK7tx8Rjd6f0oJcxSa8bzo53Bbt1OYSxeTEZMa7HUF8LvzkKWwwlOy2dSSx
gBpRBECIJOO4SC4y5ke8kdOiy2rpN5h5eM+tXjPQffz0QH/QAaXLzXiptEERl9d6
qOOdJ6zc9rIEO16NbdzUO9bY0QghnZaHh3VumsQ48gRK51tLNPf/ZVOqJl/C8uR9
umXfhj/WIex8EiNHMS+shv4ysWgvvhtH2ieKPcdv6ukk76ZukQr+sRmDju2h37gR
u93p6jtN9p+pboyU/iMGMt4xJ5oYkhHCh1L5LrFr7oIsxO3ZtRZN6cEKXMtP7I4l
tbqkDxJmGMMA2WhxY/7g+QWGm/rOwGSVXl17GrGrWdMQ8ER9YZ4qcS/c4wGIzb2+
ot0wK2y8jAo96w8ZAU5xmE2p5NrMKTHu0fwfrlG8xTVh4Il3bWIOwMbYqiQbfSD7
Xbx/V4shjelUWtVmN9Q3UoqiYBOxr/FaVVsUlLSbg4Fn9KE+KASveoY1r/0jYdzk
xTjE0rLCu5FLhwydHy6pjruP4bJ7zda8rVDYbDx2tAATH5COH/632rUghRCrZE3x
65koIGw2tfMg14cLC8xibOHDLTPa/Sw+jP/b/obBldrimoqXqZXBb5SW6AN5gw0N
9g+U6bzWldemL7vbF4Dg/8OSsCAB2vMgu9tLegVvREaKAk0cqYieQXgRMH7BHNGt
SJmOyttBUWakMxzV79xSrupIgfRFs1Adh7YTmzXriCTdyvKntHn7Xq36x9roSZZL
XzpoRE+RQ0iInV1c5W7PblezHBAEcOYsqRlfFeOpbO8rnlxPIDl9uIztV8tuR350
b/5hxW7zdkl5ccA1rYjPlgDTSfe0EolefGJOZ47YNIEZhrJMwS6KB0DgDQzZMdIr
NteCFw8D1lLFGsjlK9nATAZkegKO9XW5ePgtAg8NoikjOivuHb4dV36jGgOHOrdY
xZ89Js1q+411VCvPxPyz/2q721KE3u9WyfyigEAzlG8PVDGJwfqY5KEoEKml2TkG
tbgsMyyP7mBsQz1pNzJ1hjUm/7ekWjPu9hsMEncz7zuAm1Dw2/EV5qU+4WwYpWbB
bUo5LkkZfjcGGmBitbAwTucim4YI20iUDpjs0HTp0sO4C6kzUipfRj1fvbyDWq1k
jsRwXU/8Apd+JUh//J3hNHv1H3OyHVS6+PUcV0JgA9mIBwKb2e/uf9hW1AJb0Yo7
oyQi9v/8L5C6RIo3tISmYCUFUaTYUV6VGGLuAmtx194w5Y31MT+NNr6Towrh0UwF
Pt3mcfTLGQeHwOpwxSf3DTmcQK+B8DCLeHn8WyXMwAqA/O8kjSrlenASLEImeLWl
KGG/eso4KkyUdD1AK/BeNLin6EUNeYBBgKfSu8PXrdidA1T1RbUzzkohRXKADenF
9WkWsRQx/uB6rcVeMArkvHARxCWcekPXIBBYWaU/AWV1HhQrToAEv9xoVx0aTTwd
rfNB0WXAvLut90cDMXIWfs1xE5weamiXV/1RK6B29pXiKuIOcquRDF5kFof2dKGA
Ft6or13wp0dXIucFinwN6FDzn3ZV49I6Lqbcw8ZYX4GFboC0XVI7CJax3fndwqWE
Aic+lbx1vg2CMgcpaLCK4EsGpRCyDRczXp366RDQAvTft5ljaz9M4PTnEh2XFK1V
Yjwgbx/YxLYUuRPJsSAhqsnwkx8WnZCnkcQrcGOJ6noFtnjjE77qDCtAC2wBX/f7
rwykj5UWBqQtlBU1Aa4A7Crvg+TPuZTn2kUELE84QOgJv6Agh8pLIvYp/LWiG6yZ
/B8N3CwYMlFhYu8IMY1jATe9UdGRJH3sNO8gB40u5ShWNtGB1W5Xawv6B+yEMk8a
cLqLDR5TPLu6e3fThRtSPLofclh8aaeZ/tZ48HK28+u6z1ixNLDX7k/5NfbJUbS6
iObuN+dAPtYXvz0ggLUATyKYDXmqOSaFRAzeg81hNoED4r1bxe/OV9FtYv4eZ4kq
NVXrPrrHCdEZfJGHWo27eg==
`protect END_PROTECTED
