`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iZtBUJO/m9N5sRJWbUtghBWFfDOipwsgb3QZC55EYKSXjWOvRe5JJmjCs7qiven6
eZ49PIvdlSeh1gWgB1kdU0ynweMN0wzDc3dm3pLp3vdzIKLMKC2DQE04JEPD4cKV
gEYvyXp24FAkxksmasAFvPPV3wuTS8tSb5rxeRE9QDx9Ij+Vip8zMFIpMPpUe0Et
5Tz09gt6OoRBqkup5r2fKdHgqP9t4Sm4zWJhmr9ej8O2nmsZjNVwgYvd+1PjQTzr
u/pZDeURDcEVg9zRRraBT+bUO2TDpZf6b/8kcqqrfiKB+oQfEzLw5jYmo6zyc0ze
b7j/KxQ4TELxoMxCAhV4DkjyyrUB/m6B8M++H6DVwbF0oHM8Vvp5ryBl8MThorZv
nlm0od/ymFg3jkVLqxSUcqu26yPUEj8HcbdbOQ0ceNehx1FP3ZePYXHE9q+sBr8i
cpu83vpROPo+H4LYJdtQVl9IaYfNJJynM1cJPmm2fiP+vQx4opHGla1ow+qi7vEt
r+7EMgNOhVMkDCX7rL0pdi8ruRHHrjYfDp6dd0PPZjXp34r5mdYw1QXIqSttMG7u
Dt1yB02kC4XVo+THEsMa2/LHzbvoAjRBPDhfR00smyHEkIamHkiaYiRatB5XNN9a
GLZOAoX13hpR967AHzNmRbbSLcg0T2s0lCJ1MTvTt9zAswioP/ql78Sf+KNH+RPX
+XjzlgTIV1WhZvz6TrxDKzL90CkzBV8lqAXBYHiDm+tl5jX3Pby1K99y/Vq6a5UY
jC5VpWWd+fW/vWcz3LTcIzyPeXqUPPmXQmx+n4vaQSiWyITEjQgdRD5/rYeZECD6
NEqFLSlIe7JDnT3ky/R4OgAY3IKqglIwtPoihK875SDpDIltJ+paCnf36+6tkDfD
JQDBLL7BdRDSaG23X9E4l1FARGTZX0yuKR1PCtpVLny7uE77M673UAAzaI3L7tlN
OQB0XMftfs2N4QGAM4j2jf72NFynZ92XMFWB+1XhxBM7gpqYrT/+A0hmKqaPdhSw
p6fKys86lqDtqjvj/nDi51LMGR3IOPxZSgvS5m8d6Qx6+DfnDcCpOXYgRKXSv8xk
sl1DkqMVs1MjCTSEt1UfcJxcNT7TvXzQWeGwKhHyyZFITk2mUjHbnw1dEqHXAFpv
3Fd9LCf7or6MdUxUCcUJx4MO0yPTgUwH926tAITaEkiGxCbHm14A/M2DN0OaLXn/
O9BK6si0eIxnmHUMjIJRZNkrAB2O5M9bsl2Akn0DB8QTQFyev6gQSr+CIZLu3E7Y
PqmB8RCCkjaVm3JTIU28Cw==
`protect END_PROTECTED
