// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
LiOtram8qkjs7bzYgsa6O/QNn8VodkxLJoMVekTnw3POZTvFSPYpTpv4Zabh5Yged0lH682IgWRN
2lrp/loISqdP7MeQ1OvKZiBwMVQDcEclfTxCT2U1AU7MYQGkN1taZ3/vB8YYPxGbX5oDihoHptFX
K1skw0+N5Rtumwqz6+6GB8NunFzwy22U3K+qDFFvwNOuW2vvWHwbh682h3Gz3Vx8KpppFcjSFSsP
gmK6qlRkgn43vUlfCfwvyg+LT4PDEr9TKl8xjso69iogNgAQ8UNBRWo67aGgIpQ7ywwzC0LLuH6b
29jJN+imJKbopSnkXuciF2tnfouVbpmFfoFPpQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
0eNIUumOykX8EqSrnpRXqD58loHGh8Xl0Ygq3H0h6+UTqNSo0eaREicKK5U7iJWDqkmtFcCcpVhV
F+cqKc6KTSGH18ZeqGA4/uiDAXWLR3WooHRPLNfSBwT6J3WK5p9UbkqLn7uZB+N4uRw7LBp7cEbS
eu7hYCmZauXr60s+BI0QsRAa9yJPAO8/e+w4k5iVtGruu5PPlOsv6zbJVgtaHv+uqY833rjOxgDm
khe64dWSc9EuffPWgy3ekDx52MvqG0N8dXiQbB+DbqR/WnCLbhOiqvedEYqkH0uoQ0sd9LZVbhpN
Yh5aHpfqxMNowMc1r0QP2rzMLw6cn4wdcO7NxBBMzbPIkISf6HrqWSoz/BdJPFfAzlM6moDI7j89
B9wm5HczaZK+TOdiKrs8t9lUbyOEo7VNB4JwyvisdEJLClgjqcrYEhlkfrF40IyD4QE97ixPobYA
DYI7Is2QGlj46spBmWg4uH3jk+U1TJRP8czSmk+P50NPypk4sapiI7//hCNaPknJAr5bkjx8PGm0
QhegrdiO9iuhbRGEf6hGOXrPZPwkA4PblwrK0RLG5gE/+TnsOFwGvab030r6s9dC0RUP0UVIQIxi
+2OtQScQKXwnV4DAvk8IRG9+sx70IiiXwbQy3FbMbaPGIV+3Tn8SK8wRRMG3mWtJgHiHvfvHcpwn
SpKtBNiDHkAw58TTMBm3Pu26Lo54z02mlbFNsVNw0GpfC4s0szHsWhElvJTV8O9QdoQFjfPIYM+C
T7VyOdQPky1SuLrOFzLpPv8X+Pg4bxnIpn1nJ9eJBuK9BkHfk99HU60Jg+w8bOFun7mSj/o59Am2
m5kbLGp66f6BzNfrEbHRnJyWxBBJocuy3SKr/4vtv6ZAPMaZ74AWPlSC5m0dXNNBAbXud6LK5Fyb
I53meTVlOzs2ZjTyijsS3+23xyZhCT6uFq7IW1E+YjIybKfM4O7xacLajTr/a1zXzI5WRO+SzMJf
ZehESK7GcCZbPrZWoW5PpjfXW0yBnIN7WVfUhzQbieC/GTWGE1DrJFpXJ1Wjr5nxH8dY6dSg2gPH
1QhL17R9jea6dcUQYMyGQYDsUJRHMGQT/3JjMnGy5Q6nZ2yOe+D+pfvR6d/DiVe4VLn1hNdeDv2q
YZ5idBMhIkQqCCxYK7UVPXeJDD7XYzOHPp1Hqsl6rBronAHT7US6JUjXgc/p9g/0w1b8xHCX4lrm
HKI4hnm3TX+QXDjMAsMEoU9tYPKZgrq5hkyCN8T5gP2e9kVJCImc4IALsohG1MOB5IbuOvjKb3my
FhGa/6eNyZa9nVvgqNwuyPff8t8Z1zKyEgltIchPcedCTSVncd6tampNZRdYXJim8yURNlFKd2gw
HLLrxa/dUDcYPUQv4NWsSjn+H9M4obutIikwy3NWpo4MhDzggKJL2UxXGNO1SP5lLSU9fCuTqlU6
1lLKJLrsvjGmVkar9oxfvfG+I11voL/ApjgQryLkhnlysRPOzK5MR+f/2mURVOE7nudrh2FGwqKW
ULM17765bQJ9fqgOCXNgurskC18E7ntCYfyS+M+mtyWjAKq+Zr05ZYwnMLSyBKWW9/lo4okbURu6
isU8Lu2fzXNNgRonQFy9wvLxdvMjuTHqqig20KASjwnkiYya+c3vokA2hpcG4flkV/ziwbMya/uR
kISngCA3qk+dBeCcMfZ+sIZayoQtXPVe5sXt66nuf86oMFl/OQoahfpVoJr5+qlEsQh2PvBMOAHC
ueeTAJR5UBeETgZWD3rN4LDgmXimLiGiPkjUB6bIz9OmYcaBhZOPw5eCmlyZWXV5ui44i2G8qkfF
RJ7s8ZtuWwOg5JlLLH2zy4vvaYwkTKI46WndAavIckSb6nNzp1M7CPZbTP2WO6A54KoLAW58M/0K
X/V9NsvAkcV0x8UWKZQwNdffvfSOzblDzVx8empcuvJeKGWw3QsuTApDG6+ZTeIQ72cICVX4sF/u
1OTICSQ6oIj1AaDZR5SKf4c0VMA6bchQiixZ7Ut16UNfciEI9fDgE2D/oXFjP/vDJ6O5cVwOHjYb
Nag0MSekwhAA81zKzUUxwVYZ+lKImCGOr9hTLbqrKuD3JM745Az9htOFdOoEtYxjT38CGz4G00pH
/X3HTHIEbxRoJY1Gi8hQAIi9zzNCV845OJFvJLm3e9/98unKb6R9Ovpnj0lIylNVsLR7VPUAl+Qp
QKNMdYTNgJ6pGvW/4RGXIBA/rVO3XJTVtj1R2UFkNrNEZPmy20YPSSvfO4z+i49TPf19QSdmmTCe
y7L6RrwrkIUXL2VzYNy+OzvEnp8PA7thSBk3mT0f5eCW8lVWnA43KelgDS766cSxEFk25Jc095TS
c5R2rf/4fV1ELiVkmD8DAAMXlOhZHFPlzI3iauoKFF/I3DvHiEKT7oszUOSiwapMLy0IvlAFzUZj
f0kFAtnr4AuGV1SSSreiKxIpbKxv1nkekQQ04vD6ABNk56z6fbH1DBQLaJUdf49rTO8lTj+dz3W/
NjAqBLtuKdbQw5r9F0D0lAgg7wl25YYHIaFJjhH2qcG9YF3vvzAuAYNBBdjDm7EsUhbVxs6y3qhU
1g1uftiivyIeJwesS1U8bUQebhAASH8cy7U7mw0O1tCV7M4iyAb28KgSJNoIy5rFhsxLPU/QtlDu
IqCo4OY4xQr6WABLtyZf2kIc5AWFCF5tw3h4f46mdCraEjTG/gy+1X19vD/pkKcQCUVkQj8YqvNG
j3joXwMBvZS/ufisSv2Zm80qb6+R2lX2UByjPSafrCfXR1nc4y+0r/H63UDaL9sKYoHc1o7b6y5o
ih9r6nQHL1+W5rlUmaa/d79KY3zV0F0+AdCAROMilkoo7E+F1ODutUnZI9HNGXdwkT84qEuzWExg
xXWqELkXyZokP2FMzLMSyuAen4QOuq7A4X6PkouJX3ZYGhu5UaSxmnNjgvrW4tek4YtzxAHe4Gl4
fL3qvJ62R89+yroaLLmndC0guFcxx6wQyyCA+9qC1EuCIfySaLgrhpNo3a13m/u3q5I6cqwnl1tg
fjgCiObJKYdUY9CHKTO0NNNTdxoJy9Kqe+vSxCL9OyGZEqlLa6Hqfpd4r115M9F3SlqwHR5HmKX/
KYoVVFKJ2uFO84ubozRVfydc5GFql09n3nxucTRaypzOcBQYX85AKWjVi6yxOVNpeCSU+G2IAkxU
MNeR7oZnVTcibvcMIUB2QX5DsIoWUuW7uCsWN5EzgIZAkuwLC16o83DqNpH24ESGcdb1xiDRytAj
9nY4CqOd397q3UkDlc3jZ8tpWnIIn0D6638yYCGSR52Kz84qo/KbQyHfAcMMHkfnBg60BRMHXV8Z
6przCA43HzP3F2eBplqzenmRMiI9e/i+wtKHE0ZW0eWsVwTOfwL6K94ydAnSRQk6TPyf8CF55oZk
jIFzLP/HB3zlbte7Dybh9cjBlgFkNnITb+CGjj6EhFk4lT8xiYMS4Ar40JIcV3mhERgpNmOQdvaS
WZhusll+bCx+laC78mijy2HBXhQm3Tf9mh9q0FHGNa2dyAcYRVTYEp5QDCQyOsW4FKN8pbrHsg6b
lwvfZi4FnxYMSB9TY+0ZiD7cPJKnWJqQuUmiIh36RfZKrdgyWbyqcG4wLow5dBev2z2JtKlLXqXw
T5U59vD3gMe3R/CauvtP5ArV1SL3yyOMmasaYip9Gm+XWgdpy/+5Zt40a82AGXRWTFDOiyTYnpYd
vdq+uewI4L+Zpeu9Si+wsvTajGzwGo3O8r45vuHIRXnDKDMqkk/G+jp5E4c5CyUoY1S0yQoZEmMc
v6kUU9b1H1nH0XMuCMaPMYY6qBcdQW+vPQBdnRKq7I+SRnNguP0ZisQ7QublDIxp/q8BkFQ1W4AO
LcqCOd9fwC3cx4NAWO6JZ+IAigEuG9wjVm851Jy8EXraNt0XUP2uPno4dxXO3UgO1kNekzu6caDb
NSKkMOYTntlIdkUTIk8Gge7p9nyaLbr7mopP+7P3+zrXkUYwDoOubO7WQyhC3NbvlfxRoHnsi0IK
R8ZmVTzWUb4L5tZWgoPjhOCqJ2266PPmwGcFnql/uXs8xobUalkZjTeuPcrIfuhYcm97zOjniaGe
NVfmkZh3YFWR5IHD7kf5KBWb6MzhxE81miJWTZIbprtyuhyqQGbqmOSZL3FtPej4H2S+YO4q4+KW
Rd6AxzSgKYAZLqhy4U4LoaNwaUpeBsGXgdXETG7jcaG9XlR5dBHNHEiHkS8m0At7P7zBx99QnuVt
jpK7kDsQNGtvLIV7XYwqmqUysmA5MvMTE5LIcBvSccTcYn9N7WakSYBwA+Pfeb0PPT9fQBxKvjEa
Uj47Bhjp+KTFUkcmnmjMUpzCAmMGrduJ27CvLh4RMVXeOclzuw3sMOjUbGcsdSLlqAlvVGfUOL8R
bkiAexSKUC87TRZ2tybZbNG+HYFabtGFpjSKNvGnCRvPLtNtqJp8F+rEI4BXUNt+I2uUb+zNzkgW
0PyoQWxEQ7wRDAnHbOZxBN0qfaghVBHFZTTDerN9ZL967OJchpJUUDiRoMJbtVrsKWFiRXtw0ydS
9pK0XTZZPGPnB+vOYC/CtHiFCnWlgX88WboU0+y7U/elrm0MlWTBJBTWDnnjQEL51WwdK6gReLkQ
Nc8Hhu7/drqeqI+yr2pcz7bNlfT/S/M4b2Qlr26gWf9PyrssvV3DBYnmVeSZiNMrLTNpdWDmM7Mq
bAObkgysE04kkciJKaNBScerplS01jejUabHcbOJCNCx2LCwTcNxS1drHaZisx+R7NowjFtN6gIu
lE6lwIoJrKBCd4neLKkUwjV5d+1qxpxlbmPv2rSKiJTlWse9d7f8sZtHtMQfnVGMXYnKmxJZ1RnI
qx6uaXJpEGIpvLDQMkMUH6+PE3NTPuhCFP78vDs8PIL/lKXE0INjKurMGpg++PDhPyyagIKwaIj8
TMql1It+KOu5BXI7vDbhnKiCpZY4WYaEfMfGjkQHvCEybPda86sNWa2kmLr/py8VmXnKHMy0+qtP
ldGWvoz40uGkouktIUF/sj4XOtMZNGrlp2QJ4w8xv9e5hF2vYrMTFrcUBqyKHhR4GwBhqmTEiVmy
wm5aKxzIfwJPx5jUs1OLB9C6k7QK+CNiprAm62zEvGC5NILSCcVYyqBQSeLaI2W1ME8Nxn/s9brS
YHf1Whrhtp7VV1bQMkT0LCBCp8qvjXtJGXbF/CfyX0m+chHhnEfN4EZGBIDUcO3fzbPzfIDkNufx
7ubJdEzAd2zXhaXd5eEnQ5Y9Uv7tGHLt+T2TZGcF7BHI85T6F4utkC9SBsNTJJi0oJwEf6xiAc+U
oRVckLxjZRMQDb4oPSEBdmTlrANRFf+DNsBfI3XJItZO0uzQI+UBjI31gmxb/YIlBCSz1E4/rXFr
ENxoTTo6t4o2NevecAVPK7uJ3U6Btspi4WxAbxr1w/uJRXVxPOfkTfZPUsme83+lBckudnpxejSK
GdTE1n/KxDiwffUFk9GW21XoeZ9VLjgALI/7YvmRA+yoEyKVYIirXbHIGkdbz2s1fj92Lp97uiPT
9D4ETqxBk1cTg5sooYYo9y6AHzioISewgxp7MIA2z8nlFT7DecyNHZmrBH4q3R4KLh0lDAJ6KRaz
RkggTY+8riCVdUtcYjBL8T3jPF0p2jLBiI5eQWKi7G1Cv1RKh/K6Sb9aFf/zPvQi2U7p68qPy9HL
3v4BGEOL+1WHeJBIO9uaPkw6IZuwJsysV9vVeAZcqzsr0IvSM2WQF9LhOS1CH6nvXprNdei0MeDK
sJJTUhKv0GZn/7D0lBNzWN5Vj1ut1qVUW6uOaGNTrhikEozTomGtZGQpkOCUQuAKrle8w0wx5cRl
jpB/gfFsTv/hgwT5EGDhNWqeS5bwP6oXyjywW2wo7dElA7KRwlioCOqskxKYTNwhcwXVW5VEkJsl
FL/YZvffUuf8fy9kBIqr1Dzf+ZxEv0puIBRpfV/4+Jp9H500WlHcbAyuIxV2wXTHYiQ2j/HRk2jP
2ml5GT12kXDECcPMBjLSZxAulwIpl+7kb6nbEaehzxLD2v8UvnndAS+t3u/9EiyLut6hUvkkucx0
eXMgX99f/tgEtQAooWb9Z/UGeLb5hMTuSrvKCpLfRWOlPtQzFHmKrpW4tb04UxV1JZ8W5AWoc9Jx
BEn69d6kZxEgNt+pz1u7l+4WNXXkbwEgs0Npz7nkj2L+4W8XlESq914sEpaeXcxV1bIcIOupA4Yx
Je1jHSoxrhodhmLo9vatzN0x5HkSlAZzIUaZMzFeFq3PO6MumtgvDn49LPCFFeyAOUeMFBGSle7y
o0qYAtItnjHvWZEHrAEPOzh6EA+Hhy2NLxVV36nMndT6v+AL0YjX3VKxwTj2Ch5gtODRvEXV5zZx
cqaMJ5i99Pm/TtnU3YppDpKSuldeZPsiJG7L6xRtrYsaqdu4THFZDHXJb4lvmnoc+4ErvKKT+6hK
owm8FIcU1fhNvYbZaQ1R4SHUxYDXvDupxM5GdC7UqOYyFbDBipvIZbq6MNysZ5LF1G0lRg88ezz/
nftrzMRlw+rCISImQckH0Tw9l9BOrAZRbG/5pYp05HkgMT6g3wVbjZFxAdiru7u2sdmQbmqXKnFD
7XlX6skLmBwzAO4PE9RhDBc/aV3lF8Tyd0d2FvEKCt5t69Jb6Ix3ddEe1A2PcjqB7ClQeX4csdWl
XU6T8DK1jLeUrrRTdVXhfNFRcBVzSMKqyROzeudOJa8lr2X1joBP91negCIHfljNmRF5ZR1GzH/N
15TxAbS13ldCHBW7t0Uh7GngRSfVZIxELwgOToD0ftV4lA4TJ6wKTyj1qKIInzZANvILGMgV1nA5
riEzPguJ9RyhfFsL2zgzHmDwABzLpl+qGhpJYLBU71ulryU8hT3jsJRulG2NSzi9XEeFeRZ5zKcc
QT+bXA+u2msZuIWg6A84fGQyDQpbOkaHpfZ74YNUOxqeJXfdnFxvP8z2jMMn5FkGRfD7h2kFO+11
zFONIEoDMaGvrpa33K2HFGWt4uE=
`pragma protect end_protected
