`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bF2mpKPwrPpEYYh2AjOtttP8q0Q0Z3XeogffjklxT/oYiNnz0HufFKendX9VOUbM
k4Ups+wJlmB5dlnypPZcAKXsokpK2ojjSTbl1yEGbV4l+DVOMhwEuvj1O5irp+J5
Uiz9pdgWXRgNLDy+VJlCwXl0pGK/wmWIQS7g0Dh2a1+Iu/qcRMaDBV0c3FlAHTVt
Ec97A0QattR8oE9dy2ki7HvgBc6hmds7U6twstjFez8nX8+KqqqZ678/U6exDAKS
Q+pzyR1DkjgVOdcJeR8RCzu82OGxEqT7ZyzpIFTLOEnZ45cj4hpKq3ZCBygapinC
RXAfJR227668QxfX42N5q6MwI3GlCm+NlGrTglxgUXA8GxVD0a2cWf9qA9298qFX
7STirQqLnSw+7VnF/SSeA6CJtW/MOv8gndYXomfcSGWeICTson02fb9Kr1D/RrW0
qtS1/PtQec7KJjO5IDk3kpLVJbGhdBjt/1UWbjeJuUxLx8P2B30TUAEcucXSIHxS
jsoM//QbWJyKTPzK41InveS/hiakowFwJvnDsu91UcHIInwhCp7IXio1fvdD7cfX
qQYdPZt2F5nsvtTtwUMChbhWdll4Wy7AT8gkY4TqoqmU5d47mBmfSnNkmwUqnkyp
WnUCoj6CA1TkTDzZMbimyyNkalrl66SuLm5ZXlVPtba6HMyc40QUYs3bPhRnhROL
vaCujs91Axb2wT3maWcyoZWO7MC8T5mIrivOX0HGhNQsMlb8vD0oJQAU8r8ebvsY
3nT3+KP3VHek5qMeRTA9dgRnL3/FiO62xE+zvyF09fEUGjtXolbM+AX0cAt4ciFE
JwfyOE5aeyjRFenMJxVeMJ69ngaCM9LVV2GnyHkVXxWlAIjmbeoZZrHuySv/Z1iB
h2xgevbv12eu+Or/aRjkmOm6gIwGGnBA6S3BcFkMAhMcdLIP+G96lhTUS6EOVjhY
3872fFpP+PZtFf80H0gcXr22yaw3RR7LALaTIOQdh/ZLEEuOazoRssOuU3SPqHAe
8xsayf0TiOTUbz5MLPX6qrCOj7nB/1QwvSKlOrIYBMuHsC+MMav6gVxxvUCCwDMr
id4zyykyylR+8ICSNl1dmaeg3RnNDObbhogtH5fCoQrX6K0b2EsyQ3LoEjfR6WiY
mcioSlOfKkOs1zxMeoFwbmQwiO5EmLWdJoPKl6PuPzmztMUlLsYXPVGtunt5Av4j
ybzbP62UGZThg3a35UT53EKmlMGDiGWocV0JtqoPlXQabXwABm7o/UHJIDfkUY+S
50m5WBHWTl8ZUKdhY6Ewqh6FRG6Jd2pAcJoPyQcm501VzifeiZryJTJV4MvPlMdp
pUgv38CzlGFn+lnV5ccwvVhr7hJQXqsK2pfbUG7wx6MZPRT6Stj1Mirz65NsmQKJ
wIdMng6jP4ctRzk8yEiD+Eg7hm7YxY+bis6lfV1aBb5Tj7tU34W2epgV6RkKPSI5
6GiPWfhTuL6F6b5ZH0UoSTQe7EgzxaQB4GXoSAS80zdw7wx6W0frRd1wvEu7fVnU
5K48fot6CNmp/8YiphyavaT4UDUy+ByOm45nQFW3SwNHCHTECZgxQ0Be28VX2oAI
SVTZ32RZ0c5ScR0SlCBM4YzOOnYRokaNOKDHa0NalhA=
`protect END_PROTECTED
