`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5NNPljqIIzoUFScWHdKDS2u1GLeFOnOHJ8Em5TEot9e+6YRVL+xrrby6RUvQrmr
B+Z8FI1VYshiYz8/BhtvkvIoCVr+EXybAjJ6DQ8fBY/stTxZdVaSkPRTfwKAeiU4
+Yxh1QuJCBtyyWNDNm79xZeMWTjp+w6to0UccCg3pZdIcnhWEd5QYm6BKy6/t3Wc
6wv1N0xfdimTlNuIjiy2gtbryax6hiJIrZoAvVLjeCHEfzMJWC6hSU7vy8BmtLcF
R5nxumROCmRX9kV6P9mjA9FpWAtUO9+1zyit0IsxA+6ILBTMgmW2fIWYOzwr7orA
7gYegIiQDC6nOgfgDJ6w5lElUAMnZhGiPcbDLnuW67PJNsI1havXIisNgZY24pn0
yvETRs/rB2EXgalVscELs4BglxFruq4CSRygfKkjrHqu/gZSJluLqprQ9NUC9hhg
WtP4SvtwaLPuxfZmjnjEXz5qc6CPjcu306xYlPfPsAYJvz7CvneRJ39CKmLLfMtb
eFp0x2LJSAk21T8DDNDx9jDVofc24lkoGmMcLgxcfYIXMPqxKbO1px7PlRZyZxWl
lt8IVzV0zcb4OATfSXD1zp+RSnUpRqCmRr1RKmKLPWCu8xxluTwdYkqa4g2X7B3M
i+KlLB2hLPfzgENutkMmmd2kBHVsHs2esg7IRLB/7kQfEim7C341cGjFnVxSIICG
JLiNNp20brP9GsiQgfH7Uwr6Rdn5yUTBUrUEom1tr1hBVH6aK5XiaTsGNvuXH7E0
7C8QtRjmWJT0mo4JtDJUt+uss0bPI/qItn7PjyB1GCY5nG0dtprQ9WnKK65cF8Kf
M6RXJu8rNFkdNdqs5Doy3SixOYCUaDILfR3qYg0wAxHyqM1MrX78OnaM9iOolXDJ
tirpH6FpPfORASFBSBvDCSBMeLh8isNFuNM3YOvt0s+96eDlf1A+J/gvdtC9x9Ph
HuQmRZXVzHBp4yXcIv4rW36BaR9DGJwfSW7B4ALf+aXEHbvxgnupHr0al14lBLxx
YJaqUe8TYduoQ6PFZzSYIRmlaRSs9FLRcCG2rf2CFefwy8DDqtZTdWqFNcYYQ6up
OUgFuYybwNuDGQWqb4c8ymH44xbSLobRaBzN6iRyZY+9YefFoJiYxODqUGrfs8hf
J1zZXZJEYLv5ihLDiwbFTYMZLxRumXEMjQRimxqUiina4HLJQsD89sAGhF4GO1TC
tQD1vpkyYVeRLcl5Kq+AE8zXQUxLEGwy6e8DXNV7dDHwXSyucpHhR3SpTx7GRGMo
VaDRPfy4LSMDYUO/N6HyVrwHJ2DrCTG7vYXQLGiXka7HNvckyciWVCaEn/MF7COn
2l6ke0gVnbtXEmD+TeOsM2dRApIXb3fu2Sq41E5XGfQEiIZQEQtQJUtQrHAgkwSS
lktymFN46EC4Zk8G5yZ1IoM0mDDs2Ut30Tj3d11XhQmKXL13jbpeCXGFhz/EcMK/
IzfDkokwxlz7KhEmYID5iX8qVDjjcrTVIJsxBV3OW9xI2qIsMuBwx3ZorazRC3hT
Gb3sQDCiqiYpn04tbSJUk49stnvDtV/mQWrTDj1z1NNct+G66BvkoLs+wuGjpt0C
mSX3y+uqztV1Hw4/fTkgHdcHe6Y7QqheQelYBtQgNRJx+YlCgw4snciRdSFvi6/q
qOdBDuV6TGUas3lG/H2SKaSQEGXK6MJ/Mrvp8++ka8HWVVNx91EAWmnry2xVqqao
qAUNKBUEIvqBZbgTnF9q+gd+bxxp8L/uNV6NNiKdBPqDfEn6Zj6/VeWAre37Kipx
CL410CcoAP/CkuQSLEMSqqqNFQJ0RBPv57Rfuwq4+T005/ZqyCyJ4/tghUst+Rgq
BCBcNOllIwEYY/MnLxrtotNoT9dxPQQ1bvNaQNdAmENqxXf8dT2XYiVqERsEnik7
GurXSedPqglBkBVbgwMHLW5yzwlPupYu8VJY5gOS2soGjNM0YL4eEbIuRVHlighU
KY4BTx8goBhV1HjtY7zrhhiaJ5VFDDEH3+XF1l07SWxI5cuK91OIN+N1XSnNy4+A
oDzD6Sdx4GOVUtJVNYlLrvDm3ISa0wcQ7AC7Namv+9xtLaUUTfQWdpZzNPiTemAT
8wYfKbiTPMCBCheypT4tj1ACmmlJiO1hw6LtKVrfjgAl/Tkmdl9UEXm1lJkdfzYA
/8PxFnlGYq/JJFMAffDB/fRNwHo2i5Lt5bqMAvkh0mWuCmtN46TO1DVuPly5V7H8
2hu815hn9KGEiCnM2vGVD/iMSeK9oIGnnxhYkq9m0+F7rMflOXx7a4Jhw/3DqEbm
/n8jULSy4PGAsAwaNHQczhRSx5dE37MQ/HU02HUlOIaMMxQGYhWEeHS4iTsI/mkJ
nAMtkgFYw+bcS5mZRjFZcdlPq6MGcNPOayx/5X8wY/SVwHCnM/Tmttw3ka7W0SW0
7ueRE/eA9SPi7r+5XN2wrCGaLxoZHtZbS2MobdtYQpntQaTTubSw3OIHr1R/Jngd
1YDejARvopMdOAv7Gd9jjZIva9v9VtU8Qy5sVOJE26lPswhliRFgu96YISgsDOQP
y6If8baRcz64E2ag2Qkt76uIADLi7bd7rXkweF2zvA/Mqyt+SdLwaeagKAr8nAm6
Bo8TuAcWSiQAoTztWYlJaIvgx1Z6XbqHwEMvN8pKmWHn8+U+M1sVdu4glmafAdMu
vJz+jonYKco1UhO49if/rMwy1lrNlic39nTAQQJF++Tw0wGkPzo9SlgZ/vvPepaH
8lwzPrIIadJTXddtU/XJRyZN8ywmPGOczpE+vIds7NMxddaLRI5msiE5MkqUDBFo
tfk7106nOJRJk5/YfrMlIV3CWPsEMk+eJyXUqMBDTqdqtur5sNzfoiZoZBl8JUAh
EAimRIiLUgAGzdUN3I+SJk6nnpJ+iAPOBYV+7kQB0+BN86pGPVgOUh9Ti6/kFBUC
YKxncCNpv8Mu7suZQ9deZVOg9kXZztxy6puMZWxcr53a59vgGjskq2s8/tLAaq6J
nLu2hiKfB6XLIpEAiBphAKh5+yIZlt4CaILqNZt0rgWLf/ibOE8a3cb6lJtikB//
TY1wpmHqqAjpxV2nTHGJjt4SLG1Vd9/7DCvLm2fsJ/eYRyMsdf4uykSk2udhKrtl
4gYBfT4RA+OW5KxL27Rt4n2PDCejoxHEhrzOLg3JvxV3AlxNuhyLY3+qWr66wPsn
X4GiXEUoE+rOwhWJwd9TEkWGDhCrzZgWNZeEyPE4k81xgdv3IGSQm/YG5yJ9vmzI
dOhFEf+TwnaMp2PM4nwlOJUqlVFVBsIhbK+l4CRDIyM=
`protect END_PROTECTED
