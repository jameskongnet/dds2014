`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MkQ0eXlYJcA9dHm+6olKtYYUHq5eJeyD3rymcq5CYA21LjUlmbunOnwPfpludVRj
2mkEJy6QsPXbq9eTDUNI924Gc409oW/HsqI+iUZxYPVqEnh30znEyJVJE7UEpTS4
Gp9aT6otPuYYFaWpG0z11DgLpcGtobAPhtfHNjgWNb4qEL1WQjiR8KDDOUlUkcCY
Da9X0HO83Jq9EpqK00XBNJO7lce9jSoIvicSytfv0eafqCP4stzfZDw+c7UmkrR/
Z825nzMzVzf2gsFr0ofjBmjpnw8FglxHYxI5VxvIRx+R4r0Y9K58MbpiG2GPR7Lh
lhnTgrFvhHXVt3lQsO2SHmoiYBvfjonHagafzgWomoCUTDjVOXCH1e/D5BYBbVOB
ZYllGqv6oISgEnXoRW+JucK/qToiC8wJVrhUj7PSUGIkZsEG2qjZ7HkbKWgyi9+0
UbxfXmdZ8BQWwSPjurfMlOZ14aZgmTJFv5fJrNhezAgMGxHNHK+Xi5gBWdKmO5LN
Qm6oJ/klZqjRP08dIH99Rv3od5k3f9boVTs/Q+WNjUJrVsVqfkzSP+FSsO4lmSq/
ur/GtkEpL9UdEriESkaYQeX3sR1kSUV/cdAuUlo/8vQrnkTuJ0XckHWFpaDQFz7P
cqXFgfxNNcZFSxlGHEW0/1G0ZbwmwofPGRU0UfqPhQJ5WwSKXAaSTE6ivI88ahLW
euOJsXYty2Z7e+ymhVUGuXkIXSjzNQIijAR85n9/9NpAkOGmIyK4s3fhJA4W5BxG
Ssv6tPHGkrwzAStwndDhNhzT4EALvoVoaT9jujjERhHGJo45cIr7cmOMd3jNgWrt
YMMjpDp7pWb+0AfXYh+waBpwkiTswhZK7oxakFU8iWY9uVPntCdpfaKX+z3O6ZVv
vYv+7ospf6ocbrQ89gO7xhD4aVLX6MVeqRIFR058gBn66Im6LweD+itKowgB5LpL
6/nZbjpwVdWHYGtjtKc8lHw+ZxgJ6WT6k6v8BDQHHoHvEAWf/1pg+ogOBE5xs5+d
aSXH7IELxztYQNrpnxWyLSJSQhkC1feeJdu1N6VELdEmEhOWt1aHjtFA2VbBCSWv
B7XnFPUbBbjlaEMpMMZhBlMiTwmDvsBkUhhom6QdM6ZvQPLYmo/g5Anw1xtL3yPr
pUzrO/Ui9AgMAqqbsuJJgwK8uPQqqDa/0xT4FIFcsXKq05NKTLSg3KRJLJR6CErT
tdrnzBgRx50wOo5YFfQbjrsym+D+11fxEbfBp6gROVaVpR2ZLlOZYotzR0TFw9hT
SDHZaySZ1+dAG4OWC9rpALjDnsH34gHZo3GEQSsji7OSo529Cx5svF/jyIb1ILed
lhnLt0dOnjxvaUn4I5wrP/xdIO7+FnQlMj/ePCBKGuvoAe/r6bWCifB8W6EsD83Z
FengC32Vf2Yq6w9qCLbyFVV9X8j1mOVWHtFmxcAp0olL726z95ZDFxcWyqCuy+Wk
/lGPB+DbIVmdQYvwIREHQ2ZTkhHcz7LHSIBz5t2E1J3W6hRuh93C+hY6EXn4x1SL
mq819dYEBy1j3S3XmYKD5J2+seXSSh/Y4Mu2n4yY/QFpvtEUDkdqNu1XvE4KCkHM
1d8BY+WVYpS2fwd8wyfF/Tz7S83WVSjbLH5fa+62wC7LUxkjDPUv0EAkrbWEXUBg
f8NS+39sBlY2lJsKlDIK35VyyaXmiQ9D0V4PE1Q/wpHcKfDfPZfCOBIaGKOf4i7T
OpTbob0gKPwSA6Z0QSCzvCgQ5iAEp87sY0jJYeKSdUZ+clF3whSoQ2/6ccifNKhB
LrPpFcbbKped0gFCziuOiWqRDd87tPXO51g54WUrOyyisrXoS6IY7Hur8cji7Pab
ALSz4qaXEQJymWb2lWRqXXxUlTLmDLafFNnkfXgux0gjAPJgYNfOaMINc53ZYiZT
V5En2+cWOLuP3xUImQuGJRYvjz81+FnVF5pEm8UTpCOk4KrnDOtMXslHgF2NBCUQ
iy8QHhEnlGQWVB1Mc8ahkdEYfxhdxrJIn6iuHq2m5lhSPZHklm8GenYbchJ9ERx2
J5jxrSvRK51aFkE853B3dsrKBCM72fHo15VC7g7BUsATLCZSvEYbI8T8khOmP0nd
jpLbs8i1CPUr8L2kIh0c4cgAk8BX4X0nHCa1H+59ZnD75qwGUYSpQWOxOx34oqW9
7FL8VROd7OPW+vJlVq0JgsRTjGVz/nSnMYH6vrsmJ2q7bJi6KfAjd+hJg1iqNc6k
ENuHCO9A8fuomy5C10V4NzVNqkX1Vogtef9evVMF+jIIzi1Dm6ZZih/3jkOvain9
8g15aDyI2zn1lINRLbBU1L0jcjV3F1OEr3S2uKSkGAVz9JSyBcwDzEACOVyyVnOM
ZFMbEVHcZsaIUUVp86KMaQYGvF16CHekZDjLTwHnzlaKBRw0FsPF3M2N51qPkYkx
QENnZmEiXPJLaLt+fMUBdJDfITMOpv5V1QzQpGVHeIddPvWDThD1LpCJZ8czuXbl
GF9C4p3BvxkzjF8cdpJQGz6In5gt8xSNH71BKkeyx+Vqk7uNC65/e3b4tFKsPwJM
3dLRklOCmG2U6qq0cyzxXfR0bOwt0PEbo7ZbZU9TAhvjfmdiR/8eCjjSQjXarpUE
u5IvdGyFWCOtyWJruzK54zGu5KxkMX05E+TJj744L5DDysp+nGbuoQFAP5e+vhX2
2nu6673y/sZlUb5Frsgxrxf80PQA+LwbwYgeACqJLVzyvlbYFfBfjTQD1soa/hsY
SwsMvr1GyVggXT1AB8b9Pri16aS3HhnEZ5kN6kPRhGO34l2dKeMFK8hDpgqgjbY0
dR/VD4PkJOZRLijGL5QSZnsaPbP6SYjsOw3++fdLJCS2zJxcH9P96nbw2dI9d7oY
/RWAhAA1H3yeK1cACRglwVM58i+MSTCOIA9LLQXqv/f2PdwctEY7IPg8HJ2vg6S3
oHiS3PcBXA66T0NETcXMAsSTh1gv3V7b79+CwBAWwWaVw9ONUsPQaElvbe94fkJ2
50UWNAczOMFL9ods9aIsQIyZd8oVT9NjBfci9n0ALAkZlaKz+Ui/A2fklaotffNC
ZcguUXOnOApqsTuso5AE8vRdkifEv3ybQUG+WfX/nEQ=
`protect END_PROTECTED
