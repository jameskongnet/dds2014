`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xwB5DkSCihB+/0AC+KX3+HyIQ/jTncjxfBn1QinaFA4mLSHrwk4re/R1ZdLCEbuM
oUkSAJLwjErBWyX0p1FXh3422DbuSruizFwQwEFd0aZKNHcMC2S4T90ofmlCAznX
dO4aNTs0IR1ld3r6gDctOoEaV6DM1pEP/SXRmFH0T3rra/AQTuI4b9SqGj0zwbnl
xqEb7Mdf7iiBJdHbp9jF6rLNS0ShBpEENYB433noivvfBNvOmSteuVdkqYfs7LdQ
y+VvNbVluqo4sWtPgDETzBBybi2dQDgtwbYVs5bxBrFyOdvIUvIKONE8fxhssQUI
Q7fma/AnED5/Lf6/88+6WRwWBGxpgtn0f6IIrfLePgM4J4UvCgWJB5MFpM1nXorx
jqW7ZUsgxeZqYHk6d7xhenLX0M7V+lcUS6UutCAFc0CupQYYY/xFCDOxsbGRpCvn
K8v78F1ecgq1P9MiK3D1pU0IUwDybbGd9TKpp40YR2S7tqBARHuPNt6FgtgwdF3d
qC4fhzIi5I4YwmDxwEn1CwW9TAOy/9thc2EyS1dM0HFJxWIRYEa6o2VfzG2K+SRJ
mkwy4s3RjeT9jw9nJqc81NFMZlVsz3dcg9TpZuUpUU4dV8jcPmCb01wk/k8BSwaH
aOk/gRn0nvWmVTzVA5bJertpqIsuAoN4ClmEDqvzqt6jRKB0m1ojeTgWXJSfVfbo
RXLOp4x6dd1nQXcnva/rt2XKDyENr6m+FjX4cQ8vZ4pCeKSmY6f5tfWzrm1ObJaK
WKag7ESMvQyphUjfmAUKZ+xX4I31Tf7+3JH8xd+dggRnu15cgVHHkWSen/xEJ5v2
/BehUrOAmkvXvD17ioqHEbdqa+YxjHzd56WoN8Hf94MwKz+dwyIjHOn2YknUDpD5
jsdY+g/ah2UBV4fTkulPYxAd0+FZ1Z2RE18fjekpJmKxKo/11P3tAmHNMlt9GiGB
hwgUziNSc+wrPTRBpIO93C5WzWH4BewVO6dSny/fQb6CPOxukw8jUx9wxIQjqx6d
nS6rvsl2bpCBiOSC748SpiHMkWAFbz/GbRz9Ckr6hoMUED1VgxTZX+qGk/xDv8Un
ARJLIHNP5PC7B3XWHWHeDraOroBuRkKUFjKlcDiG4rZVoDBBA0/SOGV9cQemuAEh
dWAexOnSnVkKep6xc1bDIBJFrGp6rRrU1Z0ln70+arSDL7TMsPkcRW7XOk6d/ZUE
RiLJn8OTMfTceFbghpQS3OmUjvWzHV3Lhu/TsaegzucGo/9MfKD/Ek+oAA/cEQTg
KHZ4ZtfdV8wkfD8nr0g8DLcfRwWfaEstfIJVEleSYh43f6I2kmIlP9qu7Uut4sra
zUXsqJLmaF/mtb//Ey3u8mSW2Run6CRED4DGbNJrDrNzC7HfbYlVe5WkRMHd8bVP
KgxF6UzpNSnBKS5Xudn3dRrsaS29ZqoreAwTQilXrb8/FrYAt2/pStkfuSaGPNIr
SVvvbcHqqZl/Zw6NZYrmo01QOYe030M2dc8w45OXZqWi7YH6EEKhFEC/emrXQSfO
4tiZz70Ca/TyrLt+TpO1m1Lsbr5FKb6fyMxKDFZQw61io8LM6v8upoWNPpOjnA5m
n1O0yJzxEhyK+kTsxTS+uvb33q3/sMSAL0Xkd/8Af/G74a7JJbgqdFa+u5TtcA1Q
0QbK8uooPyWWfvmY+DRG3VVwi6nFVuGY5Aw74Ltx42+uMpDe6CMpK9PofvdKa06O
rj5j1M1zyRfqBdWbTaVGtRbwStcVcQtXQY6D/gufX8sfBTWDtyADSEhi3uJYMrx8
1WArjCFX+ADFGJWF3Oh3bnGeiZKJKQsK2Ll++KYvHHDx0TbBxds0IgDyyDhEPEzu
U7ocDV/bf9rE+ZlmxkJeT4XmeAJcxRrYSJUcRHZY28v1Gg0cWZhJ3zUiB0/BVMDV
ARdCKCAQVEv0+eUcKyROZzpp0mdS0pEwkSJ9UIJYLkRkztEfyxt0cPHtCQeaS4GE
RiOabXZMuAypKOPUmt4zcMrShq441udMEMqS8eOURRZzF5KS0RpMd61xfngh9tia
s6pG/2dWTSJ348c4oj/NE+cW0s4zyXMKSp8O6sruMK5bCEezBRbuX0rryIkkOyrl
b0w98I5q5BFv5sFxC1EbGxGq6wMbpuhYRRHFzs8IzBACxmsJUm3kj4EG2Fquqy1x
XIajw3IHQ56+YvuAG25h/o9bBCfykHNDlP+YRlL9+sj2/YNad2VKh8KJblCcZRXG
V35FdTNe8OtnK0HA9GfahXvUQXr2K0QVDGiyqXl3yYxCwe4hHS3kQ71hCYIU8g5U
uDa+Uw0/SoVBx6K0zx1uXCwwcfjd9l1yPaWrnoV+0UPvdnxNIsz6q0Xt/OaHL8PL
2gV0Mb4aZk7RzioBMdrQkdUbopqtTjQZpDDoJeuZL/PTHuDT2R0TokEDd5Gm+pc3
zQPWzp312ipVMvWhIQK+zS3x55UlYqPFLb0LHNfW99Jlw03PJDw4c/uu/oQnuHBA
9CQOzbSB0DONo9uHnf3y2n05NP/FTlKsEnDZq1NKQn0yiN4AZv0mYIkEIa/sw2Sr
o9UemssWhcoi6kLNIfpgSEYNyq5QLbWhbowlPJK7tQA4/q8pxyBbvzd+hFzkL5++
S+2qc4YV4qUQl0tvHQHcbaxB/Xvpdhps/Jv+ZisKSDPyyoN/RH/D1VxaDt/pCIo0
ayMyLqH30ZmXVqXoxnWRVllHgQru+FHdEM8uFv8lH7kNGkx5lC3UQnCouDBsIsk5
Ie1RTus/CWAT7l+I6yeaN8kzTnzxQjyWxj9ZfEU2lhV7oWu2UipyHQSYKoF0zcIe
NjuhwHdTzsODrhnsX3C7w2qZxAJFu5Br+Sn/dFK8qDIbWJjU5XrJpEx+m0/t+h5S
njJfmDKUVYffuO3FX66C/sBuIc0spsfvkTxN7a4DRoNRQ+s7Mv/tfQf18GwjqXs8
i3JkH3Q9ND+6r1V7dC4u6nIy0/dUBgcwyczZwaBTtaZVme1cqvj1YLkM543juie3
C08nV1yZd2ybDkEK56zUHUO2UOwocbb6kl3swakXSelTcNNtVisfbcEUL9Q6+7cQ
cDzz+n92a+WYVhlBquVZ5w4G9jhU2mpkUqoPS/It2s1j/Yv4J/wVsN7yg323ltrY
iZkCgMeC6FhILqcIe1KVKyXtWwnJA9k48vyNAIfPl6nMt7jJHrcuGDLhcFw4suGg
bCFnq6T20pCIlMKXPj6PQ/UFxqvvvZHu4XP8ASoQU8N2mIlBV/Q7Ez8XSaEL56Vv
BWK/ksLP83BoXSNtspmedq5Lnmn0iPzke6HZDxZLIiig1n7gx/MDjXTSibTu1ntC
RQ1+Sgr3WH8ua5dixX8AC49wQt+UB3DjWs2nRHzqLrRIkWSK4LbOVpc2IgmfShhf
SqdsJfjCQfj7qYbZSoky2wTJHyQFtAIkfb8Ju1SDExjH4Fs73Qv3vK1oye1fh5+N
H9Jixjomg1Qer5aa0HqDPdGkRK/gqlYR87ZrFvVSOIJ9E1JG/DoPSLuOLpuvO0JP
F/CxcrZCTCHqtzFXvNnStc7lavuH9L7k/SWvHajmk03uRJB96G9gzREUL8ht6DdV
qB+Nit5wtdCO3jqPPpCS9plCEdO5nlJp1f5LymNpwMU01McNQe6L2sDecEHd+eeb
b5FxFkMJtNiX5Or1ED4DbE3GKnXOjCp+yYgM04UHpB8Zn4AVvWo+Hc+Vgf/A2YbA
KkNYwjYnVqvxhqIklSPSXB0p1mOTIFfEbxexp/ZwVoXegmBUQZ3Fro6mTZPG4RSR
Res3NCAVXw6Lasi4RpGHmFaPKWuMTAQ/F8dQZUEjBDilVbSweR2+XYxARH2OGsj8
u5mF44tkKB6zdLcixFO0R/FbQCjMwbqNfWHt6dgv76yzpBKtIZ1hPlOcMQVWKcUk
EMG23nphK5ZWSPYXej+2EJP2WRx1cOd3T/scOLhslMYDNbK0VAUZk5UqRokxmsps
HyDsstsuRkUHe5iGwIsOr3HbcX+MBn3GSMTaTYJUMi1iBrZS8OnPdcAXDUxO0tjf
wJpDbj1zF1sFZnrNht4WqJ+h7Yvh7Scgww1B+pYdWw+f9rwJOOP0KibsuJnv8wQh
/4zCr9Z92A79SG/6shLSco7AL7v+13ezRe+qjV5Y87pD8qyhBQ5+yMD+AEfViV+0
FmQLXZS4454sotJbLTKHtPYUpTU7jxFYZAz0dt3GLSP8Ck/5izX1UXiqp4OLH59t
nNPdcDzT4mFdvLvfmO3pTZE4+3N8h24QPlNHXXaDC47DA5ajQCi45h9O12YI/sbJ
umjwX/Hydtc3I6/EaC4JEJYL9oXdspqclfiLnB1AuDFBYbVzMEuqU+f+JkTqUdyb
K2ePFhR9nlyQi3oWBWhNpp9MTbHtyk5yeJFn5hVb5Y45FtYMKu/3a1ICpO3KdNX7
9b27wD/FsuoOHvJua3rBNTsP+je4weFBQNDculA3J6hNxJKQnNjVgb4Ot2E8xkuv
FRcd81dTdwq8zxM/c90gTKRsriAWZYO3udPRAT9oJHcqXuhHADoDiov/ZcK6eSWt
WrEW8hET7F8WR9ExdaZGlIiUuc6tqzmVs4IF+6onBNE1h8ogSzCACa/AX/1lPC+4
ZX2zod6IdxMYxAnlmqGi2WJ+Zz9p8YxooYTXJXnA6qSjgMKuVnL5dfo2C7J5ILaG
bXbtS04H1bQdq3+t2j0EOhXHl1G/KaaxiHUQLfKcr1lpQ2mfdS9bWVLlDspyhmbk
8h2fvfe6OsiwIfYlmfytyOrWywCjVkwBD6ZuMztk5hffMB/8MrF3nhOFZGEmZUdL
SL5O31QByIWGX6HHlzei8/N8/79ZJtHbuDWSH9piv+GtWmMyUMNyQud3Aj30PISl
5ZA+J7tFGGWav19jjip8mcdRo7rYFvefsqZGel9hD8bwdh1qssKz1jIDWvmUdq6t
U2RiPI50cjRuG/5a/UEQREhzci90Rx6034TcOyBj4T+/WTx0kYssqjqfqiIDSU9f
MtpMl4C3Ad5w5+/uwauAGzeYcwvJuYQ3KL7lxF/009CZWeAj/loDy4ASHBZM9z0m
iQ1nfEUOqIifUrtO74T4NGX/4l0i+ovpIJS8ApZncC6YvrEqBtx0P8NVH1jaM+vb
2uIDOdZazduDVby4/wIpgYYOqWYjSBhsaLWu0aYT1RfPAJtXO/zo4IJfu4rr8Nwf
sED/vtNiHW4KVLXVLcXqek18eP/SlQHauLAYSkQ1VVNqFyJfObDdiCnxLF2EBjzy
Ov5GqAYBn2ITNdEd683A6fdBv/L9NHqEAbEdUmSCokLqAmASqUDKtlrJ2sLOO5LJ
M4JD4wpTt/umIkYFCfqrRMVqoqhrwis43oGiJuxePfiQCUORJaWL2wkcG1JWr63P
uV9QtV6yMZDef2ZKrZe6LJY7Myz3m6w/lu96abV0srITshfeP7Pcvd+YXD5lrllm
idScQ9pJBUq9sQimrgRdoVB/1Yhtc/KzkG5z2OopvSyPaCn0MYtAp5nZkhx3sCuP
Hl1OU5folyybs4/Zmv/NyLCLZhE/H9yeh0xFboH+H5KZJHbb3iNPWToqc5DKBD/t
1+gAv7T5Yu0PtOB0qHFkYI5d9GFDK/OfbGgvAFD8OWkfKQsVfBSZBZRX5pu0UiaK
+HNQUIka1TDr1hiyNjIiobladLueQ+oJbXArrIcQ+nN3t62SKjgayo7PXUFF4N4Y
JwrecWbKzT2MJmKzgEa3MQyF+2ORxioZ1sntEYM05ZCEPVAc3qY+NjjpXPtU9qXf
6aMQdG5rF8TS/I8yEMnYTTu1QgrK2wjp82iixX9Xe7uzfFnwR3Sz9NFOFyWmtAqe
kyY2KS1Bjkx7EgDqRM2Bou+PKtoKWRs3daP/dpBHYu1V2ma8IlpMYK4D+E352fUK
ST81XqDvBEvhX0Mlg1iEmOGFOH7cFCgVMD1BCvIxiwncT6vegTmYzlFLChyIZWL0
5uBKSMmL+AbyXSTq7Sm/7F8AYiK9gMm7Ihw4P/03svVcjoSJYpqPK1jQjw5og8Z6
DRqR78OdaXJUYA5wpINUrJg7xxwAg6l8b4HznfyFWUaG+J22a4O801tCKITezUvB
mH9Osm+p3Y5uZTTYVbMujbHQnQZKfN4Q/jTn5slcJprisuKa9O7nVfD/N9U2qIjI
p4gj7TK66xFJ1nK6P20gsfLCX+Dl97p9fPM8MaXNzlS29p1VCzbdxX8+wgBRo2Zx
HquhSEUKZEUr1ULW8gii932BlSAP4TcOYdQJTLl5Oroyug3kqxzLQ8vNCkPD0kRN
FQWQeecBex4WQBj/ObovmYlGKelAHSP11O9Mr/uiKL8aXVbl8wEOpk0tIci7oWfX
82gcV+f2BZVxrw+SLaGRAp3Sb+ZV6RVu8h2nm3Ii2OQtDjlEs4DZUC9Q18P8xGxQ
UfnV7lLRezCNAnscK5KPX1aW43ZZtsDkUkqn9eAXINF+CiK6njhrVOkdHDl9O6Cm
9VfU0mnWQRgU/aKvAsaNLCTP5BGwx620/bR8xE5B3576BPfoQFuyrpv3gmyM663M
Uo45PQR5tKRPcDXNpJVtQFZyEAEegkLlYsQKQQTLQMQ3TZt+XVf8TRrXJgYo7VaQ
8Th/2+uasEfR7xSmNTU98VRlNO1kYL/itf2+ZznCwipM4ArLiJ5iCNastKq6hQun
p8cJkeTk+Jadzjk9y8KR+ZHcfRL6v2G0FvodFyUCvXj3YwO5liyTHeT+WXeYcrQv
QN9L2WVStzyt4GyvKxqdHlhTvXA2tMUbLEkx/FuRxjiCWKR4aK7KpwfFsk9KSoZw
wlnrYU9lXnr2LWFqQhmNYYPxJ26GzL6h8Z1kJj4JbxZuF/+/5QygGJdCOFAebklz
lLT8KHkz96VPucq14S+38Xbog9bhQmzZvmRJ38YSpEzwByOoQaAtKXffhMBTmP1e
7XeT32ABaoGYNMvX5XXFLfVDRVe1+KyBBzjUY3qswP6o+6FhVasu+zRbL0Fzbs3e
bkaFJ4fFC8Rz1s3FpqODfvCbzBb9q2dkPK5tSrqgSvt6MxZnFb65vhg77vPBt7Yc
DZ2s83FYjgoHzj0NoiFwrMen/oiAeaqCgPGPHS1vob7rCEnGQA2nvgg9agVWNaWl
SBN3wDlTc3ZB3B23D9WpDqlJA3OIIKThFGafRrerc+AtNZ0zWyRSf7+7KdcwShPS
vyr3Lo+eTOp/2mf3hZMIbEfs4azwYkcacbhcyeKCBaBIJUn63UhNYIQH/UffO1BZ
a7den2kkWoOcQnmlwQOC8NnyHXoItzkQ6nSv/oOM5cB6LX+MrfBbQQgBb167xuEG
nDJiyuAnoGLiVQG2VijEgFnPQe0h72PrpG4wMYSSBkjAI4szk2OV6VN5a1IRMmE1
XJGmxFUAx4q7o16eNR+l6ur0K5fBM2U0FHQuM84RbOGYB0kCHOHWVLPp8jheumQ3
xqbJctxwpK65UfAsUMoDcnJlnm/0D8C73fzfInRBzfIoP13/SFjZrCgPD2VYfWXf
2XLPu6xospyT05VjyIaWAMO0qDUDxaIWfzdwo0TVZY09scsl9mz8k9c6J4ZhSMmO
qnwHQ7r5MPYJjvrLSPGZM32Kr2nYfq6PfUvuCWfuiCqI1A65gjbI1Wi/u4ZTUH8J
/16EzAsJL4DACnUFS5QNfyfT2k96qSJujLp4SAAZFyZ/LkxYMaUcBdPQWA0tvV+b
UKrAP8zpfiFsbeBzbJ+WY2/H/QMxOYr6fZsTgJ2Oz6d/IhboA0nEXRHydQlS+uBA
aKOejhro4a5wR6EXbSYSkW1fYNlF6ZYgXwWxKkrDLt8ZXmnhY0sZA8zyUAaA6OAa
6PUauHpJHggBnhRpvXGASyPbQd8iX7beKJIz3UXvndqt+od0AbBUIED89AMGPVzL
/EEz4LW0yFDnE6A9wEI+Qdhjb9VU/onSkG9SVy+syUMeJfebYb/oatHH0vAChQ2t
71u8wuToT13DuxoiZKkejktXS0sS7kqsDk0ApvPUrOlWADcpDjMxfbHrBnhTtJc5
2rodRHm/gXBy3eIaocmCUPEu0ETvFA+75QjiSiUpe3NRTq2tM47NAJJVV+miWZ+3
JmR+rUW2jak97pWevZ55Dv7Z2D8xPLq5rU74kpDij6pZh7XegJpXOwfglTb/gmW4
0sEN+YoRPF0cQbbeKPp4BckXY8gkN+wdrE/4qBa4Jc1jMLcb9XY8DODtziX2wFgx
j3kTOj+VIv8GlJ8+PrauL8Uw+jRagGnFvWq8zhFP23vx/4lmWEpA4YUL1HbbvO/L
jUsciwxwWnywVJgKYThc0ip7Gx2A/k6ov180moehFvcZUxiz/mi5pJ1N8VBWNo46
et16UQIi4Z7FSsX002Mgm8JFqBerKc5o6mLJ1dic6Rp3TnmY7GOuryUQboFkfkug
VNsrVfU4p70PX425TzwYlkYUmVGu1DLK2ku0wp8+WLMxyo9+5cHq8hQ12SnhE2pH
2rY1KUkPhBUtemPeWK3ok8Jw/amCH8JWAOcckuM41SuV1R4jd5KvFl1+03z7tnEo
Blvd3gO3LeeDMlnfik4Ve3ITei5k5zMh1qA86eVuSm4OcgdegdnejBAZghsyyNKV
mC7mlrN4uRqXYtzCxjhocnKxcVKnlEh245x/R7y7t05ye6tSEywMe5+usqFOeV1y
fjoVN4q+nt/mrGGRJKveGWyJS4YqPm5X+drK2LorB5voaLUbBx0wYPSZdVwdKy1m
iGRw3S2vLfn1BLJvChEd5221W9/YT6FQ37ruHldktJDXbH0eLQ27f3ikdQhGxSCK
wjuYvZlW2sb9Ly8FcRGwqAtHmLjDC7ssBVGuGFJ8nquu08IQPkcAdWboFP+v/PMr
cT8J+d7vvN8zxkXw6B2mHTa+F8N0FPT90rQuANOEODjpYidKWqNONPrLDVks6Yly
cLTtcx1gKqZ6azXB4xSXEczscHpeOa74lVY3RNxjQn1vvBwpdHFvZprkhDM6vBDv
1YsHHUETVgjGUjGPkVcfOSYc7DyBDPO3mSeBANS7EWxeV8CK0NS9rnzJh/PXac3Q
rqKv6hTho2XcigGwsVOw6sxyoAQdxmEZPwPQ0YL8tlJSqXfY8pO/CF2c1hSKMx9p
MVK164zIRRlxk3nVVGlt0/+LAXxL8yvK3J+fBNcEU573s+wE6HG/roYOiWPGffJc
0TV5vCD3GixfY2+tzOHLQzif03i+RZbXW0IkHjbHjFlpo6BNMwL9XVWfdpkUVWMK
SAzJ1rdvEGhThYPRfJfG6nRKvMXK32qGDYXi94nHu/8s9u5sZU72DlZehpWt49ri
wSZnz+rJKJKdMts8zAosWUgWzOz8QLpyu7e/DhzlsGPoMimCXhtoVyJ8dXuo8RaA
almY2Bc6dbhXi2r9eHS1cUJMZ67IQIDGt3T/jvlxitJby9ZCZfV/NRpNtYzCC8H/
V7jIyjMdNKq3qUI/QPNhS5qUCzkp0LEZsD7762E6pkdhj6Y9AfhXlN6udJTOlblN
Ou1UqEQecSk02O7/Kotd/crY0qpP+VhYHHYTuWErYhn1sQ9i+DWH1AwNo5HtVPWj
+MA2niinQWESLoILQQAqDk6/24wuaYqK4yZd3v6695PTgy4/g3dCenihxZmn8W7f
eGXPLFiNOjQERdnXEPa5lOr1WHY96dDsjlrNxbCBclS5Bh9ehyWR8frJ1bbHbYA5
FJQHix4aHY9sfzwAkB9FOVBOoA67T4JLPGcYnxat/UISFC/KGwq1BewKFamBTwkf
+3mc8lVAVsKbis3KD9+8xmk4VclC3I3ME0ACbjtgeWhWMchd8GRPXTvsp/Z9MQme
lk/CEJd/GAiyAPJ8NLuL+p450dd6QAXglp/wHeQj7BwDAL3IJX1p1/uUCKrvWXY1
lF38we+rOjLlPBijZgi/L+WvSgCdFx+6+iQVy3SLzvhWx4tvn1ZTqocaHhJc0reK
Q6o9BKw4ZLaCNoB+D4dgUAWeRaZXyQLBqwrUez8QBzQrnDv38QJXQ8cy4qAsoFMn
OA07ACmb0C8tGth+GwrtXYBwYR2xeWnu40krRGGotkgqVfPrJjNSOxEfbh4+vefg
zUUfRPFpb+caWiQ5L+pYmcj0Ezg6BNGnn2HFx82AOwcLYV1/YcoPy5PSvAB/xXAO
mBcUmZPka8fW81j2GzOwuLWHgVBRymraz4C1Po4tNV3zA/Fm6irlCvsonnq4cPt5
x0DF7LRmSJDqBlIugSCZGf9GDbdU07b/VJcH91eHPyGFzSSEVY5U/EupQHu49st6
P1mI7pQ1bdSFNiW47uibuSyTc2yYiDtWxsck63WTlKgjV1NBlT2g4uPISrmFnAVl
EB24/fN6PBvVpHMQ9DDabgU3g2+RyNkEob8vmTxrdRYLTwtjcq9JqKBg4MnQsf/E
sL8hRvCDvB0R5EK6imCd5yyPBbs/hI7/mJjxJMNX1WonLWVf1ouQQRfvRkS8//zA
ETzjYu2bimpOFHwlcq2VEdrmv8egCvO38piMWAvGPdTyPqT+5EIG4/j3Fpz9Q/yN
1aOW/65wu90OI8GIY6NFGIW32Vw8uIsmYbJzfEYc11FvVinxHN1lNl5wXFaX693b
TOuCOWbJyeI8g2sLw3kIGREWklhQYzBuG+UL8GDOpUkPftaNA1ZTtJcABCpITFsX
k7OM+neJaUq+hiI2vI0kzWDVafWh3rbh6gv8RguPl5ozXTQymRWfGzQohHfLMQ5L
D0mtTc1uUyLNMPFD4fPlZe8maBq0nVgIaXhlFB0iy/+mJse6vEUgLi8Gmgl4I7PZ
ZmlfRlZNiZ6Y/IXLcOgWaf/gXZKkvuOnBWP3bS9Qz+Y=
`protect END_PROTECTED
