`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vw7pd7usHdtODbVTiwbWjraY2preyNnhKP5zMxI6uULgOKAK7/+FDo8sPhq1lMit
N0y1aM2tLduZmcD/Qc84gBXHYJ/SBDPokVAt+AadK5ooRDY/KV98S7OW9kkFHPH4
ynvpXU8UIEkYsDuSeGfg82vM/xupiksvuscQUVapBhTRZBbStoTA3/2KuuYE3b03
HocTUoG57gZp6OamKrP0J22umTPFc+VVBLcaxCAGP027GmYlIO+sSgz+h72m7q2c
7fZB0ZPKi/CH6oVZhLOI7rtAAbZ4CvDvTULfPN06a/W5OBeJjc4pdBOmmGx+3yGg
rfNI4gxlA7AYsqPc8d7kOxmJ2J7w3hWhcrBIg+ZbBe9gO6EWkt6xSvBhDBQk1i3Y
UC8aedYBxUlWXuXxMuXmETL6ENqhjt4Y/MJjtdDO/T5iPUlrUoapABA6nW8FK99L
a82ep7uhHNHv56KDnu9VhC+095XcMgk8dDHXk4zQyakd9ep7l7ZIullHWnnCFUkK
AMYUweb3yW1IdNtxmXjz59kZLvtxnNG8y8B9pR1pjRlc7WFJqtRrdUzxqW5OvocN
Q0/01f9l6diSJDJ+tBvuiNygBgA4QmlsigF30pM4grEc2knbmneigijX8c5uzaa5
GYpjzFBxPmNb+LuLOpIiXVWtPZfDVPhGNWHTtp1fPsmyygdig5sAOHfQnIYJEaGi
oXOLMQn+3yNwzCv9t/jtxr4OJ8zbBSF5J+PuU1E2cf4QbQCAOU+p9W2g/6u80ioM
U8EXwVUw++8xlINNvF5+ANLgZ3naYJzbOycH/7LzRsA7wPQaCRg4MxYHHNCCQ17K
hYKkrdsXLtr0OMXxJ3fbjf+l9eJTUxTEPT9nfWUu0Yx8xlF1nhLNwGqOy8CEw1x7
8/HOt8O5zaV6hZ0tpj6cYj/ivgCvD/nAzKS1Gg7JUboLFft7JjP7EZK++nvxk49n
EuG/H7uDiWlU/e5DvVJhoRMPac0b00yMztVZL+buWIDB4M90S8nBWOQCnqWQHf/A
XkiSRM7ssIdsoHr15NLU09qL4jPPR98JMXHNMdd7S8kGH2n+y+GLeMkrV2Eku3H0
+OLfGFrJGyqIcH0nAO6KfNCkHJhRT+XnMZo6RoZ679QFsAonOYwoUfRTOn7XI93f
i5H9Oij9on9bEZooH7bIbqYNTK0yJ2gyoG64S1NdTmvVKZ/Xq1pM3qYhiHJwOKQD
EV7jkbHRUPyY1rWdviFaewD2ucbEB2BuMGEfQbgZjVYlgQUsaRLmeAXMTytpgq4H
XWdTsqMyRZ8meUw0rhREf+TS4JuQgryNn9YB6c3mSAu6I347MnHtSksyeYmFltY2
WGH6lZQTNxR153lt4OU7sXyrpn3lgqyVnL7QzXNBopJPwezebAJBgxwwypZ6yIiQ
YaPu5WDUpTjE17X5kagD+L5CYm7QhfjmKq9fBxPNAhCt3ajor9x9G4/zP9eLcppv
SUvECirSQqfUWESmp3gIrGCZHM7s3ASL3mxKNh75BqPa9DAARMoRntq0LZUSxfnm
S/6RHZ4afqjxAwkg8B+VV5guv0kE6tK8YnBNMtfxXXShHe7tynY6UhaROcVXHJae
wxyjcdEKPya9GMphinvA9eYQxKdLU2qgdTA5yukMhZR4zlMoUY83icBu0LvaO6or
P7BExj+cVNZKdDYtpO7PAeh2BJawitA7gxmvMM9iKlbeYBsH77GY8bIT4RZFt4yP
5aEo8klX5Qn2UoOp47Ml1EpExDdT7LxWygX67s8IFVeQpjBv68OXyB9G2W3SfNYL
5phOlARTlkKBZL8v5OmU9Dy8JtTf9l/4mGvrjJ84sKDud9LdL146AkZCKmoj7QUG
2LrSyOKBiRcEgpv4Y/5vCbejQnhPVt8e1QstC7+2tElhlvaaGoKzqNJGA19vVHvr
`protect END_PROTECTED
