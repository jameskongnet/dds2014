`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IXumo5psuPNXNYZ8CBcGlWeq00+92Bd4vU1elVq4qfIVPrfXnsIzM6WhzcwMhlM4
PJIAunsu9K0khbU1GIuVgz6dJB6YBWRdmIuo7hYHNbAZFcPJhk32EDGJYSP6dr1q
BvgEiz20mnz7pTcypww2DE2qc5n8k5cMc+uSdXlHYfSI8rt2ugy0t2NTb+4bERlB
blcgqNN+M5pqFKCtLl50QZSjkqv7NZsEs5IvrX7tauoyfOAmGkWhI5yRVYO3kJ15
SQetZc54KefPxcKmER0OQArzISHTkTItviJleD/cMk8NPDukl2JxLotc7KCymR/g
aBkQX1pXWT1+o5BZA8iCkJKkWEvWeL7JMfdNUWr1508rdmfkUTJJMDNlw7Vz+ykZ
z7uALCgTZUuuflYXcA2N0ad6f0bCpIvj/di2d9sLr6ZbFKN++4LjNUcP97SUck9c
yCLDeT4LxaOGY7IWrPEfwZ1DPBx/Z/QuizjXSp7CXprCDJQ2NGRgss0I6yA8tiWM
KgrVeR2jlZmX1IIfOo376A5JpKq0xePpYp607XR+rkY=
`protect END_PROTECTED
