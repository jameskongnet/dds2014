`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UvZ/INiP0JJY+Q5Vyjdu+gvrjpHiEvMwMwk5SuQFnlUVtL0vl36ux4oA/cV8qnvT
97/b8rx7iWi2+2pdx3kN673i572UV308zy3Amo5Wxfc1uGkX4rVcLlABtJFSD5nU
gi8sbso1VS6PTQhwRz+esvTFodF0AdI4yjrc21KbWqPDW+NRxljHDVw/cTfcVDYZ
CAGfwGMs2pMROpjSFiBGX9WwBH43D1AXXSYqz/tkZASjR9L6kX+PO8gFa87kAnRj
KNdIzQkKoB23FIV6UjeehDjH0WVd1pyURoVNNR+9nXH/tOxo5wLnsp3vGVtPoTxB
sYvUdpdtoSNoQ0Ef3F3K3eoIOtlsqfd+jillC0UA/m1PA/7bcJUFx0FRlwEtCL3N
8Sv/TosQaufBrdOMbgKDnrIh3OduklvS95lPzjdrCKE1REeMWbBQGCW6bGix5WhJ
4N4k2OL2vI61iBvfgJxBgNxWo73Cu5S0SoFb0atbiRwEQ+r3LtfToPa5taMTX8aM
7y4BMVvKaHHGcGB61csHcyo4yp5Hxz1wzs+ZgKdWRvJyLoGb3viNaOmKJGLyTUSM
Ph8cMuMgEdguFBlgtBgyqYi7lw8gu5rbmvvzgNm6nrEk/gRJhJ4C4RypgEKHx0Gf
e9U0vRkHXLr3bbjRYMQiGOuAR5+4V/ok4Pm4yR7q2U+7kxLKufgkiniNfkBG0har
IvkE1YwtgZG6jvYAAmDr3K/aqJv/EC8a30M713l8Cyxapn+mynob4lVY9tKD+v/b
PJfxh3WWFVHYWCij3CvMPC22YiEfsiPGQj8X4I/xiwysWnkNh/6snbjpndKsHEho
4aEvxBq7nJ8sdEx92IMICcuuzNB+fY1XGgiBpw3qDuF7k+cj/SscE5PrURjPmshb
FUpmA78KRjnqnk/XULQWFwQK22IsKH2X/OThuk8ptMMPpZcoOTyVi/65jKJtw25u
TyvGuoXcYB3DoySk6gN6UaAQlIqxbrotLwJ9G4ZoQE46womGcoEeBoq2IvObMLJ/
qvD1nHwMkPyVp1uC3ACerutvaz3De4g5kTToLEYe6rBspF11Ki78O4z5efvzbLOw
AmwlLNxfRnnYPi+QNFA3J4CwC1kL1FWatVSoqPOMUoOQYvCem9hsBAD6EG1zR+59
Jt/we4TfC0PtkvWhCuuIRv2OTnlMNx8gPgFweV+mltiQfOn/KJxdi9JRQuFMiwk+
exzLQBHMhRjE2M/kQDjDHfyaTqdGJeEpJJJq/vY/71y1elthJ9WT/ohcI3LD2vCS
ypCYlj+gLE6VKi4Nd57etFBr/oXuLSHbUJ+9StuXqxA=
`protect END_PROTECTED
