`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
10tp6KpO+Waqj00/6yxOZ0q9XdevS/e40wMOTE6cjg2dKnqYpG6rnLWCZtAVaFri
L1q0af2JLahSgTWBc7lk5BwG2LExh6Jychv6gB6OGZpMGPmQeY7hjs+994kkjwgo
Y2dNQf3rsK612ObpD8Ib6XGChXViCMHGd0qtDA+67TXc6rBrsc+i9Nuz9xjKdAO6
PJXMl4Jq3r5qcx2+9AGs2cvvTlygbr9E0mq/cFJmiJmNaNjnG6HiYKzsxvgDkVRm
ha/dtk+ve4jgQn9Aaal7iODlRgGOylr72Ikijten6H3NfGbwcHkXD5C94yGUu/Bw
M4gBMHTN0Yp1Bg8LhsF2hVMUOMP/nDJY6FAHrPkDoGN5JxxK9qIztFMscjCKrmSv
/zGxtLwvwSqx93AkI7aD0Yzm03OUVOUn5XCnp5ekKExPE+cvJdzzaCbp4QKcIH/l
OB8vV+nqV39VCuoNe0PplBlKFoQ7+XWQ1JVEEGKoz3udU/ZsTNaTaReXTWcMOCQN
MEBqmJgkbzjCApNY6UNvuBYxt3S8IvAN/RwgKqrMtH3oM/sAwQJj/4HIWcSrQ324
dKevxW2hnEh3NQZ4R1pjUNiEV5RT+KP1bhtFDGkKhst+cSGiIj2N/lgfn6b6CqOw
RfJFwqtxCgUiHmex/FsD/pEeQH1TYbBnCTeWODUJ6UBxIWT7DVTQN1EX7WtfMQEm
P1YMz8hAaaH0l0wUeO30xszHUIseTX4IONQOmOKezH18aMzYM9Yruea6X+ev+N4w
2a/SNhPFyfoIjqwDpreu1cMC9yk37q+1pHr555JMaczHWJTMpJ8AI9VZy3K87TUj
vMeDKwx90qMKXfxBO1dt1qycY4jyWX6AA4TN5VuiLf6RV7e9eiXmVSp8suee8yZ/
bbXCJSVxUPVwumY1rl0mO8LS7mOLomNXwZhFXv8dtHOnHvRZkz7PkWy2nZYtVHw9
r2IP1BAh+CI6Lk+DTMgaYnmMuDQTUhK04VyLAR9cd8YXuvExUs+9OFha3IqABHWp
OGEXuzZKQafjBlyhLjk/FJyzcBbGsxDKmQyRLyPngmEU6nSnQNhlMHBAFXoCSY96
rsT53EbrYsBQ43v7Iwh2kGNbztJ3t/bJ5xzya81gbqONaNyChLRL/WWcvtIM7WxC
EVTOclJHwcazlvYY1rkVlyOS4IKZy3ONiP1V7jp7l1uvwF4416RjiyAWa2XIIgR6
bWjQ0MUwTwXUPG4NPSmk8B3dLPXsYqyWGG0OIu0F8Oytazm+M1RYsTRgvB1Y4lXB
afRvxexkpxQn/hEaRx3vNTQKVk5Kr7/h97MUd7n36UEcLm8F5fHOx0q4OYBUUEcj
yWLm4FWqXDGMRP4Zq/jmcXh6bSd9/ebemmzOmXh7+pftarnpx0rHNHaN+MmpBPFN
kSJD92EIAjBqB16WGI76MzIAnjlkE5GfRorFX/HymQgEoLv9QB3edn8+E7iWOkNE
JCB2Zp4WB1EAz20VDDvtIbS01Y7CEXXkC/9xxv27HxA6soPjfLDSWBBFU/T0MrOu
XpWCVcNPU2FIVA9RAUqZ2vfRXqJwYFbYltwUMuZQPNvMxuVgcFAPOVpFm+f163pO
IEZ9+hkEKr2bjJaNS6dEBT9KyUpFMQwEqrtqkLNVImmsR38ZG7PEdAFOAm9kZMfk
io0psZpsDr/wljr25TonC100V/od9xGBQpxybzjvNMCbOLhM2C6Q3qotdhpX5NfC
azeFvOhylwhCTIIVVPmXPEGsqtDVW1zkn7x1fclsxYPtzbMDEh3FgsE06buxSqBe
WAk12RvCxEfznaKbifCqwvSHwWm/PflpYZ7KJ1CJ7jH7leyteSgi9yFTOhCHb3hs
5M//TWR8BmJUZo6JBC4ntEM0NWZ7OECn1sR/ObcPkWbDaQ4YzbsXhQIcgdGRKBmK
oCJMlVN/ajnGz45eKCIQT9OtD7AT5hwIxi0OQjCvaSjt9kJlh7Iz3XtSf+gz5MlA
iSmJTR0Zq+ucxXoJYemmpnekmzgnYQeSLHPLl32+QdvHXQ4/AwJaD3YGQQ//fMla
TDcumgdYhv0gnBK3Vpmcx1ZlGyFsRpRmXkhFH6ZtqA2cVc+uOS6WgqauTlybc5M5
nlnqwsX+Q84cx4/429152H2GC9J/5cz0RgpFzuszRTIXwQaZa/vgaY/rZuZ0Z/yv
C063ONvgjPKrqTOxitTKe3xjVTAtBgMpuGhlIThKIj9j9Ossa403s4/47SbQajEa
S/p146oKwCTnwy2TKFXguAEn/6WAzPF1iyrvdvamODkOj7midX/hbK5sAwYlan1j
TCO+iUhihDBaB0Z7C0bwmaUxILDyyCMI2UzdvUQnffM3iv+zfWd9mkqE6gJekbcx
7fhqDTyR/M6TPQsQp5FZhSNPJAB+qssNXntH2WnLcJiqJxk5s4F6Wgna3Ry7V0DH
XKzlEOFwbEkb22q1jI81j2gQUyXQqtJv5uqWHGam24h+0ucmxtzcuXSozJzm3ZAl
YTpLool+4FXcNutfZIDOCWzHkA/bT2Fkc3yEXQtE5XMWVsisCCqXlUEG3ditbKHS
UIhHNR1E72bFvnZFVmKvCcFt38kLMV151rR5rL90ErUGrNcCB7i/jzqEo+psPGaj
hIM4ZS2cJc2EWDLMdqvIyXBjhYUDouN5Yb1f27hMzrqr900jobp8i2ya91OjPksR
fyaJqdqORdpRcHQunkUxA08Ond86N2/bUii4uyrruB4/ILjzYKfpao3+lC358P+H
/Hr9aIyOns4qE2w/Qqt0hR4TNayGHzyIMqz5+WcGtLyOAl/2O3IYaGeNzqnuZnY3
bGZeZXVwz6BZ484IZhvbdyTKJHXhjetfZ46Jo1Gdt9YdqhysDujx3w2dSQWYWlms
QfHWWwdp8VW4Jezz9JM37HWtQvVjqg9TBcoBShe0kf/HHHGW9s8JvJofDp50ulYP
NQlYgSXVrivcKr2TwtmEWNlp4Ci6YGGZJF1ige/A/iPLjv+fEUaHcMh5OSEiwca9
lVnynbCivoaFcWttvc5UDaDGCCieML2eJxSvoJPiBzZIacNrhnjS9qSENIvM+O4/
Y9ppicajX0xAB7vZ3KZDXOyVU4H5rv+AncnGK05xB4V4oQIONchHI7ekDzIS4fJN
GlrHvs0AMdleFW1aiV/WdCIfeX/Vo6hzJgL61sa2DnubGHyDwdtMERDX4YRKu4tH
f88qINiEkrJc36riuwplxs0IApcvsRwd1lD7nf1236kzqXW6q8OuL06Z/M+JD+t9
G673oxoomEQGrfW2I0dkq9T9KiIddkdfnS77Gde/YIvATYJ/sOk1bsNBu3JEhOIp
suGf8ZAsgcy+ntbN3AjUQEBjUNuCHJP/GkoxYTB0ILi1Hzk6jLBfUeonstCVy093
Lx8JQ0rA6cxNdZkqo0zeojaeip2ears3MK1loZkGv+FNKP64PsnUWYgeEGle3RWV
QARicaSNVQEVwNPaQNOiGOkMG6Qgw7P2TWcIdj6pK1JiIP8/CtF8DP4bRsac+6NU
l7y07seHIXDofT/dJbl/8TM+T9GVm6exY4UqFEvRcXoj6gZecKDUp9SUFUgskkgt
2I15PBNe6Oj6Qsn670o28A==
`protect END_PROTECTED
