`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5JSoPWPA6oXbZkBlYAsuM0ioHUKH/KLrZyHlNmbOAaZFe+CkSVCJ4J3dNumGu3qO
6fjuKsnxN4+FZ5Wwg3yijos9xtTxtQxurbMLlyJexb2VFVMC7RkpLgGMAR/7Fv1e
WO2/FFlxwb1mxd9OsvJiex0n4IH/S+dJW0J7TBkvEwvuZ3PyO3zyyRRVEboWONzr
SSUbd4x7Ml5q1BfwAF3Y6qZhfFNfFd+C+HlkCGWIcJtTpMyTzGkW+Y0pc54POaDY
10fYqqEoX5Kw6/AnapshodC67DA+QLhboyMFVQIVp6QoIWocxO4UTbAQhv23WI6k
E49Rryz8aAqk0rEB5DTTWaemZ0vM/LUOLOaHUSgZrI35xMJjR1/VoKy1F2Ymy3P/
zuoGCcNBtN/D+QDKqZw+4eMXyVQ00b6kv5wi0KwFfq0jI0r0AtVLi8lTcCZQKTwt
JvYkQtKEhNoKWv6md73M09KGdRZ1oUt2fNg6HpLwEW1vMOaIhRP9ocvzRdaHfRzE
MWiHhAT2fEh8SvJk0eIM0btk4SMh2bzSJdorunA9dc0fiyi8o34pj5MWYwF32F+P
iTiE34PBmI5dpGeV7qfFqGA1ywTfu89YbjecX6/5QTQsu4m7nzItig6El61ZbsR1
sxrJG3kV++Yeu14zxjbMDuxr8kzMvSvJhVazzUXH6nPRD7SQV0FD235948onkHHN
nDQ1z+Mfq6wR/hTvk46gsTqUbOw1VFl8SpQ0MsPvf2pp4huLxdU+l0n41XIO3POp
ElSL/9molqeLEkbbCPyiUSAXk3msejJPifTvUGWA7NE/onU8d5Bw/eD2i1VYvnxF
UxyXjcw21VYmrfyuzd4yzQ==
`protect END_PROTECTED
