`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1nVxF7ATp8QGLV4V+Chzt9OkrjgfsblxHWNGP4rXi5lrCCR48zCP+D4dxmApOZhG
xFR//kw5HEvnDEYtIGbVMpKJEM9lwWU3YufU0t8GkWe6QG8ANduA+baoROwAeQH+
UKLpOlhTr6DHlOlo+x/TJDu+TYo8YN67ZearLc6Ie/1+iFFkziho50qoKhosBvrh
mnoyfcIC1TZ23BCDPSxIz/D4aDhaiDtrrrCE2fMyht6YQ4sNu7ld01I3QwxGX6++
T9CCOQQ/F//m9gf0ubnZx+9nz0j4lcsLhmI6r5KDec097fCaM9gAk4xjKsQc9IIU
tY9EBPU2q/GBB8JINiI/uoB7mf57E8Le+GIh3ZUQD5gHMOda9F3MvB2W1t7x3SvV
+5X48wMclK5KXFG7D5qbv7llxwAkZO9g/CB1ANYME1xTMh2ZJWf68WlYGmr1kRgW
urO+dBfxa3lD+/6CNjC/TIwevyvOwq8JdTM3xzrOrGyw7yTr29+01XxSRSnqzgyB
iHVecUdRMjvxwi8BCulQ6oJSZyA/JTOw19thWuU5McVs4Ee2BgIk01SSGtsn02gD
ailXrn4lT0UNzNKucn5tYZs69lmuNM9b6FuQcoq55uxuMSW93IUddMayhzNWwo50
b3fVMcIU2cwANe4srXLhZlvpavEnUEHXGbTKrtDIgTN0fJCn1enFT6YMGhlxASE3
BgpQQ/OWrfDNwFIPCVHwU1y4lsrpU+18+mlwoLth+Hlp5vK+IOKyh3tGsKSF9r7F
TdcNXGO5+nPAg6dwpmjfcQuMc1wGFehK1CMdp3MNS3KXC2Cm5cTLXP02ukVUL+0A
FpLYUU9LrFGD9QNFsph1kGQ/dv6/+E4wvBDXa/YbNiMeXdZt2Dh2/+G0L5tvo3gW
+eCw3E1lM1kkW2Qdd60t89NAP4g4rtVZCJoN+g4PbT2J4qypx2IkrRk0IxPXXtIH
19BDpNt8N/PGWrHX11BOQSeR3Me7f+K69baQwPlVTgQIh4q/HpgjqzrWWHcug3w/
62+t3W56SVptgRPELugDHUBU0g5jcOc9vaYPjSW35/h4APy7OLzXw7X1WsKgsfaB
Fcv/hMPe7kmePj9bmX1e9zgK3v2i91A3kweiam0bzPXYSI4UGyh4csfZ6y5O5TDw
1vzhLEsB1ZnnA+mkFlzfVCgT1pRH3b3DRg0XviqmEx66GyYPUMXgYUiL4BoadRwQ
73vMMv1r3j0UGFNvHjY68SN91VRumAdVUQveDRwWW59p0f1NtnMmlIQ75PST4Nq4
slcGtdIgjAX7+TdkBs9/Msdt8k5mZ2m571/0puhSEOeI+3iR+fc11phUC7DOOYuQ
7bILFFI35T3Za8JW/R7spR+iXgKDK6j7dlmG0XtTS7risFsmNTugjoItk3GU1/KG
IgWYt7wf6ITy8FsHjarWBHDlA4nK8wGJLaiLtqlWZI89ABBP/xGxduX7OmmYizMP
MUD1GZWIIyr8Jxpk3YAwDhWqZvsMLgy1vlgqfeUmLNOIc0ymNu3nfM/RvZSreA2M
19fJe3RPeDemrv6AvRkFJZ9SdV5EFrxEhplyNW5eK3N991RRoDDRFiQMtEIm2odf
Q4IM8PrZxfBdldvnvMnbdxdlBK2hyDIf7FPA/zrqB3nWBzJjWzeWsznc6NAhqQr5
8VVgGKTN5sXJ61c5h2tr0ot6gnHsBAe08Xco5s0oD0qIoDIB9wZ3d/XeVB6tqlRA
V2BrIB2B9yu29ogEetvFUpTiIK9NKSZ0C//XP7cg1dizqS9BJEjEJCZMYOzahu1K
WjsAff+vmDfRht8V5i/zNMcXpc2J6g+AkAUDrnqlrYIWt6SsSUa70ZaRZy3EXgui
Ygkla3Dwu3HiFEpfoduyEJ96c7rzgOod8gS4wNL8om0868gugV1loJnADe/C6a5l
w9TPG6pRHM7zPt66jwdjRtb+/a4hn4YF5AOEgUUKxTkugkH3GQ7e/R8/E5j4gNr2
29wJhVJ8rzPYutl4v1kvO2UYkalVFJ1aCM6D8+8E2k8dAH1dIENB7tmdwDIQya5m
hCSjeAI9JZIZ1kVHePm6zLE0fMtummfN4Y/VSvbfC0J3cOGaXEoRDG5uXb47GTev
RXsNpsYoNHVk+QheLzV5NB+lk7iwQ2fn8puc3CyNR2MrRzncsU4c+Ew9rzv3m4dX
r4IidR76VNBlDUCfd2mSEv0AiwaBrcOj3IT/aqsV9qOnfvyiPqTWu/AhLmM7Vxeu
BEN2TZfXcG1XmOj+RDigJvVdyNKtew5quPi1b81KIvAXSpbh8lkJ2voHZreiL/SK
MulumdARMYZ4eWDGUTpVKKoE6tyX3x3QrtlHUU7SKRqB1Hf97WEJXSnFGMvpLNtE
Q6heUT7ErNo5EhR3jimM1sXll0NJ5uGerGLp+jUEf6eWe9np29Fbw/QhXimr9b6x
gU032BIRPBKhmIgkOxM7ashO7lWhKT9RgX2751CNMutroD6slUZIL+Cedor9ErZN
+lWfmuDXEl4X69hU31WvCH0J8/FFAlMVOaSaIdc2XLOW2dGa2vePMHpMc8PzCUJy
s45/hB8N7UanTIriW2BcfkzFULe/JcEqIFq+ndOF/oFGy7jdBoc55MglKfJWXaZ6
zCrXd0K7Z/pYYnzLoXgOZjHCTdTjBoZHp+YobeqYnH/c8prn+8tCVV0EyzIF/Fbi
f8RB5SDmPjdBsaCNRZM344OthBQnEynfzFNbD83raj8uIvaS+CPvdBUxZe3tv5sm
rlyuPdmVcDjEVdyusRVxM0dMzjRcUf5JsowFDFD7IIpsrLlKlTm1Klh/TqfGNVD1
xtiwuKfyX3CT7MOtpEw/pPAwPI/V1CVa8qFetuCMyJ9wOY0dKGhjjIWB/pZce3uQ
HvWq2Wnz2d+YeeaYb32W5aGDK6UvyjjWTLWIpAGpepgDbNSMPDhnxPsVD12Fur4q
XZW3Eu5dJGK4IsdzXWRgSyW8KfbT9DCktTSwyDOILDjiugmRyCnpLi7d67qDdMeB
ruzjmcoKCzzq7cPxm7+wdHoLvMMtYtWCD1RepmoLHmqdUlGeKnGpTmS5Vl3Si+Wf
eZFzsf62dmuFoqXB16z2QLZhrfXWZAALO9rHmTmse9I3zJVist5P5eXtx9FSW1JY
jWhdnFuQWCRRSVq1PWoZF7f1NlbBCH4IVRNfihpVUjieJJT1a+0ewwCIw66uuFQB
4u15F3eLHDRfK653D/2rqDJiwCkyxP96dtE9VT8GnhFR6ddlj22qQLQ4NtzI15kJ
WxcQx4EJSmlB8KSp2HEClXwFXD1ITtftdick2E2FwGvn2ApmmW17dkMiePSM5VtW
yygQXuEGBIk9r0SzhM9bHmur190ECTYp2YMZkTKiaIvITyA+31YHl591EBh2UEfc
FfxAhdvlcQG+r5j6AE6prKTL05vx0w9WLRzMdTSjhgS1VgLhwb9Nr8xhIvFXvsur
YdCo6Iz/S3mLNNB+F2+Xh4zqMg+VzLpK3HmB96ihCkHUT2+3YXgdYx3D4KJULipZ
11KvnaBPruCg2kONUkSkDJH05rIcwcTdxRw3PUWDbbo+xHoWD36EM0adFr6BTv+K
zKr1oRzxNLWbf1AXfWBxltWfbTTznGs7aosEAW53ucD2LBRTW769rekcKKKL4C2j
wxgXopFAZsOKK0qj7PLlHPLfznRWGFLcHwsOw3XTAVLgDjAFObI1kry0VV8Rpeqq
z/yssNiuUKXgu4RWHmfxAsnE/UdAqMOS3cgdpMs4p/gbF+CI4ZbxJf14GOsI/jFB
17aFEpbqM2E8YJp5sAz6VMaqlkIvMQBWRz9iBwoc3RVoTVRUDP29CwrhW0RSs8EP
iOD1mG0+xS8TWzAbiD+Q7I/NoAAzkCbl0y0A0Sd1UfKmZw38ZyNVyZIbbZ7wWZBo
xHr0LWNGtSiH8zK3WodY9q37rvQGGEWgKO6U3AY1V/bQiOE+kw8wUpGXXsv8XuFa
RrZsylBO8OMwc7CTlThq26AmjDa4JQZOz8B8VtEWJo57rnZ1o6ldyiTVZSJLfbJp
PleVbQ7bkZM5EzWW4g+115J27v3z23heKU9A9j3JvcB19BvJEOiknhPTYyEz+q6z
mAQB7AtFC4k+5orcju5+aR9MtHKB6TKvW6ceyDsaUubLDWD3F9/BWVBVK0XCTa6F
V1e2eXMMtzZorYE/ix0XGsUZmiWHv9iFizp8nihi4wXFor8xdiuzYTFhdgqF6s84
q24myhYTFDo/IVOLHGDYJXTRth0AsvRjxU7cvIWfbrTvWYqPlYhgApDmukU4Obnl
VErqXI6jAH1epo4Jx2olAkOplAhi+4h08NyHm9C1vDax8iGpKViDdW+zC3Pw3xDY
Qr63GXdyNC3n8s+dlWh7dPJT0wi9McD9CvsL+yeO+zB1HkH2bwu3FVKCQt/jGpRn
lvyWd0WHBYsYstlgQFEKOjeEkHI10CpeG1PruwCFA9vwWW1bilEzTc7uN5ami9S1
qjuooPghfb1cTuLSkzcQArmVNz2CQiUL1ZEdEJhN86cgZ4fpGX4qjEORP4r+i9lW
t+sSOi+H40e8pVIM7bEFTFg74k2eO+9BmvWTQcuLJubeOfQNDZ05eCjQOTVwXUnZ
S52ApDi56Tj+sEo1K1qxwManipJnmRyRfNOPzVG9A5W3R5Xt5jjIhkIoLadWW3lc
wa+AmIZLLSWK/MVNnrFNZYVd6krj9FX7NSaDiEIDabdhFbmztBT+e9F+35KX16kR
TJbMnPfgES+7njecLPiKBqjGqXG/dVbSawvt5lpLnidt9cAqQDwoqkrymc+xONcV
9On3ok5zLx+27kYZXSdRiGYuXeYFh4vXcCCemJ5dzShwMLWEfX38drv7EwzGm/qx
ZkR0CQKjB1Z6CATMTnz5h3GvUsuLBlsfYk+AijwUrNZFVzLNnFkqxhpYoP9vnqxu
ZtwwCgv6A50qjUomg0yAMFlehPRMNnI/wxRKW0PBrdwTEjrK8QdTqxC52ikMqgfe
EjCSXX7bYovk2Y+z3YdCVLcxtZFfq4hAFVq2UGwRdQkUS/Z4ZY50TgzTYyw9/6DJ
FcxM5dQtzTJF85tUqWUGx+1yNIs4G+GUACupnso7A4+/xfO53+RH6/WUZdLcsCMu
k2T8/Q72L/GfwDX3ReRWYKFfmKBp4RAmE6czlufgGs9+CgZzZvtrLnt+jHbMr9M2
wj5sJ1dHA+YJBeW8CqciT4cZXnDg6G5xu5Y+ixNJuFfr0qZRUFXeIWSY/+IBXi7n
E1N54X6VBNEPYiVzzpxGY/hBOk2xVfybW1UO6PXVEkgl30Ey+qcH1d2AxSpj9wAj
u/8NL94lJtjhiiXvQHd7NXWspi/81uaYqvV23AYhCm5yqkV3W+3sVGtqj+oJmBvD
JG6kfOfb/a2L04g9mVmB4OYCsJDwZfpJ+gB2GymTP2HX+8omdr4KmMwt3qZNNjLG
EWmrsijT0ftAQxFq8DGV9jKXbja6AiDTif5t8g1eIpKuecAXaXSRKvW1QXE0mGG3
w680duB19DqQNSyg8HJz1LYz7L4sWBC4N9EfNtkxEQ32BzFJU705sZgjSwYmarP/
nF8BbALL5bht0SAo6mRBImppk5JJqDHxYT9i3RozT45PjnD/l1rEn4c8XMLbtIwi
5A4Hg7kV1Ul1vPH6khDCKlLEjDTFM8i1oFUNX4/k8kyBfQf5AmHUIrGhVRJLUcGj
lAINh7lh8nfMEeO7dZoLiYcQDRPoUuNLEX90qnYmuEv5mAkdZl2gVLLMvRgJURrk
qVwulDzJXFxA74zbHSfOI87bjAfJPHHvXkcjMMk8kx9+dr8/BnRfbzeO2yDaKO2j
GHb5l7vhn1U9m1HwLvrvGid4j2wQiqKRM8gF/P0FC30jiwyThINBxRts4BOAk4PB
/zT+9iH04tz7ZE0JwtrarbfqQvmXtbL96q52eTDHa+snzzIwvyvY21Ulohf3QaP8
MnD3qxPneVro6yzVkL+kw2RRIY4/KyqLmgY8deb56k0CxYYOSn7Ebkage74Hso5U
WIr1IPfvG3lOCPXtqKi6rTHfq1dzGHxZYEDz4xf5kP+VHPNkabJSHQmFY38nBAdJ
c8vry9zh9pBQsWZotLddK0DDmnGYBMZio6Mf+WEgCIumZ862QW7L+mjWF/oW9kso
2f7A/QvmUV1Fk5T5M1s6Ld7aOInbdgLFoh/UQAxv8o11T+TRhsnwzC/r5p5Fxh8E
`protect END_PROTECTED
