`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MJp81/wDsRqbVE28e696njlwoTXL9y1wSp4y+1E8H/2YoTVL/6aheRxuJUocufls
+fP0kPcEC7MJmBkw1m0KSiVMiLlmRzirAEiM0gCTem7u39S8jybKQ8mXvN5SRcTO
T+vhp7gbuZsmoHj04GHTVSfCWFNmG4iDZsSf4G20kGXXxJNNlWe2i6SL69DI/u8Q
cMUUxMfv73Pm81tFV6j8EDjaC7xVUytWV7IOnbJsbsFo1/Yg3BDbvscpRehYfxkd
lbNjkX2XkSXyRwKxw68dggY3dk00fNKJX73tGHE3/VFKcPI9Gkc2cDp2nHE57CE3
oVJjimkzN7hN79gQMPQRKcbzK3VJndvVlXnCpa9+6hJMtG4zl5csWepQIXKcUiSH
38k0P1CQ+12pUwBonq+HVMAiYu67K9R4oL8ovBnpP1pzui3SFUVR1Nq+n/jyIhE6
UdBjxZ+xdly7LtvJD+8esyTV8V+pQ9O+fdRzA3SiyUEFbnSlSqDWsmAPXEZjU+qD
0qf9V9PgaU5McSG/Ucf1NZnbcH5edkzkfx+SSWdBMgCi62jh4DBGSPtn8ThfSeJe
b0C0osSIATa19pe2pkLLM8mPOI1YuMZSjKBVFB4KbCa/99Ph4a1O5nXcV0X15oyk
J+shuTtaFpzdpDQqGUAH1PtN1kuCN0zV+2G8moBM2VlikHuALdSZubYCpWDouQ3p
q3WJNfxF+FusUmQoE/994bTfflOuBBjsQ0bZ9/Uh8so9TSP9sgrcnqJKK6jeczJA
gjmDMwWOa9CUyeiRQ06M7YTYol/ymoo4hP0z8I16aCMc+kZaFaMvF2Lrb13eBVLB
lEDUjD95cmfPrTq0qIpXndPJYRSebvUxPmqbN/Ux6Rgasw+MlHBDcddCV0fFcXjT
80SxujykSvSuEacG4CASMbWeHhDREzubcCf7LP0y83oc+tEkmKs+JW6TUcjcLf5l
UbIreygW7nTeRO6iW0eNMYvwGKaRPGhR1UHJx6biphIT2/Gyuj2O3ThcgHMtBwxO
2Phj0mjZxsFsPhJuNP0q9RJOR1uqacaqiUNuSPjBVRf0gecjZYHaetCYXfgbr/FZ
cHatVgTgdf/LrUGeARdhZrXCbxjHXm9vl5+DptqzowfmUW8LCaXPr+3viKykaV8t
Xi0mBsv9m1Gadka7KJJWgScNalBjeg3+F8EyEEtRPt9zT9RX2oypsXm20f4uzFN6
QGXBQiymuLDlk8NXDdR/sJmwzyBVSTLoNeRxQYDNj2PkIRlb/fm6CuD5QVco/fAS
4f+Rn+5Y/8kDnLDLtJmCZ0+f0pVN5hv2v4FjnzG6HEfcgvOfodAAfuaHnZzgVPFy
5mj1QwFuLN0EZGGZ7GR07frSuMI0DQMIK2Z5VaS1iv0NQqfueOiHYv+KjgxNvXCU
HqqgtziuBvujc9N3ntN1s+pWFZ/8cPsnbV73NrjyU+CRrAASgxzWR1gZ6Q/yEBgO
eeZNJQIg7k68yJlQVPzrKAAXb1a/XvTGbrSuAEbd4IkFyIj0uLLzu8mfeu4iVLtd
ZRNtwtDcxKyetB5adpL86YPDn+P5BxcoSua5SoBoCTjWz867kqNE2bAFaw+DYw7J
2JmnG5iqDYy0gBgf7LldiMvgAubIWOO0ceDF/QogTwQcdY61fwe/EZLsmde4mW3Q
7C78uUEnprz3HmMGPLdgPxX/wdmPHVG0PgwielssGiNkPo55xgGi5DKlrk1sN+mZ
yoPeHP0g4zX/F3vDiM3VyWb9qNUDIBu2V1NB1YejLQOe+tzSRVRFuBKdAJzoSqBN
KQ4NfgyQBn2HgFBehntouFFv4IwOFyhHfTNHfRW+CtTFw4XVdv2WATOHjG+O9/8y
1fHp1FxM6FHkeQJftVkjgnw5QeXy6Qgg/QhOhLUhpcdkBRAGR1Nmh3nMZIthDywo
Jr4g4vKVdHs8gmDuWpgjlITrXnjOIIYKhrRxYu4hW2nBWQtlNy5rvUDvKTSMZn+u
F1Kf53Z7ama1fDi2ms+ietaxBTRQt2uoRMkt7O1jhRhndZPaNyuklmDEOqnCnBPP
W3FWK93/SIlvSJyXEUbDQiFC9MgfwxxnAbra9nYBaX+Mnr0g/i/4sP0c+sC0c6H4
tqAV7eh5E1KacXAMYlNvnQwqrBwV69mPwG8yCZ7pP/jq1m26lgtj0kCMiO6SBrCq
9LV+219oRRPXsnzoiT0Y8NeUZ9bYDN20JFf7LXPQd1s9k4atRWgiGSdUNH0gCJ9G
O2LT0aWhXZRyIpD+OQ1aUiAGfJLSH/ZOHYEpiB44w3ARb8zPSUB5ih1+o0q3V56r
0ExV1hEsklCXj1X27KnVcs8l7ufz0ON4lA3BseqQEJXpTopWnQeoG08RPftnGmHc
7K1SIlwlIoOalqygxLGD8I3ExyvA4oILP0AX9COAnaRXF977SJDaDB2B1477i3LP
yOSU4indq0OoQWhHw+n4C7qnnY/lCBYdeVo6CEBHsHheBVSF72tTug/BvFg9yrda
tAWuqSiKwEli/fD9jjk9FpgyZTj0uK4rfrMLwUYwzYRUGM/sNJaI5EW6wyMmphox
r6V8HUIgYFdZwY2jXCGJ8G0S8aNGB6G+LylnNHlvdBFXgzHKTs5qP8/yE8V4iBsz
+ac12rCtmHWM/Be56vo+5mYKCsEf4ojqteC44JTLxAG3Bx8ItSoRrpuwK3ScX5Il
DNnbg/cWXxKHaOOx+o27dN52OwrvD+BNGMYApfaLxKxT4kl/jzR8Xi/bTjzHBWcy
RscLXoknwOPVl+w2E+Ye7Ch76W9naNHOhmt2QUQvSmpirFKHeUrFE2yqf7FgPAYf
CQLXufPCiqWyQllVcjcTpHcyWlPeJhLwQeVDKnCqnNphNrYH19CSjl3oXdG5EEkk
odm74p14nPSiRx4vcVQa8EVd3SfhmLhiZr7wCxjNELagW/VykqZDJP/ud+4GyOoe
OoIU/B5Bm+ycW2t6IEkIehNTWy4oGa92AHPAdqWjdEfLQ+wU8FtpsE7xIHFzj4mZ
qxwxtjHZCIhZyxnGx0MOeM5CU/xAiA+CpjKraZw/ZrWITtJD1XMr03j21RgeFWnG
lf7tnYXNkPOVXSmdQ9+sY/BOh5Z0ejXbMxBymyAAZfY8O3XR7jN7zpwP3BnxijZo
qJUG4MqDI0EMYBhrArzitxCKjMqErvNEE1ic0L5bwHu4UJHd84jl59H2dP6MZJi8
/rtKPKaJsrtb2zkfm/yCpy2aNz7EGtuzGM2eKCzihuV4A1fxOxFzraQAoSfFSXT1
h+DrJrb7/d3gh9NE2lMnpcrt8SqGpS6cy19VDSYyUkV+cLMGda0VdAoS7LHqtD9W
s5U9rBuyOF2Xt0zsD2TvojtRQhCR2nJ7QCkLFb3W6dQHJU0yzKiczevfnXCQF87s
GuVjTpXyBOj4ipcploLu1vPd9q7KFNQP8V+iJphLlWhw4DR4gD4Nb9wu+j//IRpQ
T0eVfml7otvrjVp6FeQZ51enZpJd3SCVeO3WTyhKiH7cxZ3dawS0VKI6nNmHZ464
aiqeHzkgUi31HN+te1VasWmdA5voVjins1G1aowufLsQscao3ih4W8mz6wxiKdbb
xh6lRh1C6LLtkmw1BEWM3RjitTLaolHSlHQUEElpKeBEgPfOGpQSql+yixJ92E4j
by6kD6eIHEPiQjosNM2chrgWLbiTjeqQf0T2ZVL45DxO++ypnbhpWa2Jopsi1NyF
mgZF5Psv/PDadeEVkGzXvsnYfAZ/gZ2GDoi08/fAQ86/LYc/KTP5K+vnZ5aniib5
EUNasQONIaQwKlOUIynO8lPOwD9t82bSmaS6tTdYCXgWKHf8V28oPmHD0kxNMNSl
/L+x9fsKywlXcZ2DnkmHWXHz8tN9Vi2r8G/VWqvBGl3BfWxLO69RyUYhIkRL94E+
i7zBoxo0DQrgzSdmyIJ5ZtqyxdU5Fo4CmmApcOqv2f29eBA5iAC3p9rQFhIVy8b2
/Xl9fCYnAddGcZFiAKWnuqSQPT9Cif+qKXZC2yUzYdUaBr+W9cNUDDsr19qHcYP1
0HZg6+c5utGI1gMeDRwMI8ru6e877mx+McwLBDRinhGD2ioTS8ZXRrNhEJ4CpfVa
`protect END_PROTECTED
