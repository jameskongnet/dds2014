`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ZkUl0UIK+/s6zQqUFsCcvJF+EV9Gokflyvk+1yvfusj9IAeZdm+3cSvU+5zJg0r
U7c3rOb4IWQDYI7GV3EhS55lLpGoQH45AVnQsWCx1XgGmk3FrIcJQUrTO+5gUUhR
i1ImuMP8d1M7noVixgIV/q+W7CycND23pMN+p7GqryNpByGmtNC3MGAFdRaAub06
xIImYnuU7vJ/JTpHHRuxt53dIdvzhTjaJwJXfJfAXy/SWfG4iwJTHUjYfFC2jXU7
1b2Mv4Jut+B9Cma4LPn3OqRVOgBwt5siO8jwdk4YDc9ecQHI2hIN68gBCiS4w+4v
h8lsFpFwDdUErYirM+u22PqKtFjcsTLaaUI86lYhLppwzyJHcNXpCrcupbA+vGS0
8JO4uNroUX/gFWYpjgAh7WZoBwdJNZ60QiiyKOMhhX9Fy1bDRCDYXMClCXMLOdFJ
YCJhQpHoSHBo+nL7kdDpYmH5oe/Bpe60K5a80RsmCl3zdJ2ffEDcw/fsV4DxWg9j
GycSgQWjlH0s6Y7bmjIKdZz93q/UDf5/rasxkVYdkHUs43f9N3XjWuqG281hb+Ys
B2TFgnlRvhrHa+XEk4PvCOgHqiK8FfKWPbsTa0M8Qm9ud9uUAPeg8duuhhR4PUbd
wxIl2PVOYubNEX/1uBQQSQyEy5G6o7wwzAEggnW4gmcZpK1ocKv1ICAv5/gxF54c
e1ER1ScgzLa3pKDRF7F+jzxEHVpzkWUmDjPV4tDhjIJ/2uSLIqcXaTuGxhMG1BHM
baLrgPl/G9hRF0XLBiDuL/DkjhycNEv19t9YteveKgZWIRMeFH4syHEKy0AFUq7R
V621syDl+Lzrn/ai/XAwnR/qUKlAYjlfCgnT35bz/RjmTxiLvUv6AZ+70TbzuITR
1rGusXbjF635E3bKfQACi/Mu9Les3cmkTuHvO4y++7V7v/8Tq2ZlabRWe4cGR1pR
2A4XoYvx04MWfpSa31uVT9JM3oLeZpHe3s592vaeCisfcqI7GlCEmRCLZfkWMErN
S74yi2N9fJKBLzHZfwGpbtmpeu+1VnhkDKZq7KR6GCem0sWlrcxAwM/WYbh3N/PM
CrV/FLrJ69ygWfxbG4hFPYH27ZS8DzFhx+J5JvZIUecunVJtlCW/z/G6XPNwi4F+
i3xFJFXSFCynwOJmnPp2P4jFQ2XQlBZ+zBzlKTN/RZkFuZl2gO5GMHtFUL6STl7D
GgVtW+zm0jFKw9ZuOFX+sANmTiodZBE65/w40p7kVaKDBy3aAJTN3NgC1qI4Brl9
HtqOOMBBTyeaZ3FwSmR//cTBgSGgzXAM2ucv223qAzE=
`protect END_PROTECTED
