`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gUmNN6pqrl00NmfNpV6vXUoBLK52qTHqpA/wIh0nxREJH33QTOjOFPnBx8NUZV34
Tzk2ADPAOtiYJft2iQLTcaeMIbsSGmHTH5TMx1hg2puw3mCjZRc+p8W6kyCtRRDR
kP/nkRaCZA3Op7eC6mFEtWbdISSsC8IrXrOQgl68imBc98TTNkKpKyhOquQjuKfx
zWMGrkYSEQkf3sXEnw7NxrHj8VLUIUSB2Zv/yOl4OJMXNtj6kwW3rEopYuwj/YCT
RC+oQsqjJrB+g/jhLjzrpQeU8+aftdR6Tcwqi4E0M72Bb1D2ZuTMzPPCv6tW9/Z2
bwWDFYwybuVl6Wt6uQn6ZOeCx5tbG4SEHvFeoZz+WQ1zFCeMZDQfz8fVB7Jicavh
8ocylTVy75kwlV6P5+FGl+wP0m0WP8vtuulmD9tV/P6g2cPyQzB1Ps4IA7i9ae13
muyxg6BSDdzJKfpgFZwKYSMciWoWyiltKkleQkTH8m97uDtAsVbTsZ8Utj2Lb/iO
qfQpPA+8QQ0YnimWT+PtQ1nFCtVKZHbFAb3eBo4Das+FKxY77A6f8nWhT91yyzSs
q7UtUiXccFS47hHEgRJXAkgoahqES7/m38zeBJumG9lQ99yBFO65Q0wV52kjA+Os
9VSlW/SVf5rOfqBZkC213JytU1p5jK5cbK+YKicusK17/5FcqDzKI14u3f/IU0gQ
GI1ASTE/a76bAOZZU2aFVi073YTSeF8/IAxQtCYfyRQBQ9UhcJGn2xrOPWWD+3R+
ebaFUiuU53uRMs2MOP9qSihspQdmaueTyiyUMFGdQBGuQ1P9gO3C8Uro41th5zbL
8TLcjn1UlbqSTRemBXV0D3AwjjdS5R96dOIOmb+1gFn9tV3cL1nXuuyNljGciP29
bHLnFC7vvXrCpKJ9CnuSQqi3Vm3QeQQhupiGuvu7tQerk67LjpSIH5R6G+u9ldqD
iSY9YORHybZKFhS1DwriqiP1sOgCZazvUFrtL3UCCGDhwrjhAfr4Dk/9csTGtfmw
oWkvciFCn650l4zI48pQniCvFOFR7Did5KCvb+7X0OryOyGF2rlNlMyw8ctpBmkr
emlXtfOGxPI20m/7C2377x3e1/Gw/l3zGwZQYv26ZKBQcyD+bmSWCDDLZJIMaph3
EVej82FXfzBXCXQJ42jkvNwcGiyB3m4cUFrs0kJ+VUBIHhFNYLs8bJLRZzgJ4pH4
r6VpvDxkn/FlmT0I7gs1dl+oxg7mbdZfh92jbD3Jy+Ubsiq9YbiQqvyIqchQ1Bal
kcFOc/Tct99erN3NtrKRCqeMJSEf6TAKl3T4G2TcHQKB1gkVSskQpO/8hd7NnAx3
XHSiwYm1e6Gz0uEUW/IqaYjUuTo2IokNjDsb+yS0lesAAaOnIcb+diP7dYd7n8uZ
BzrBEZ0EXC3hffZVHQSXeKrIaj97oOLhk6X/aJQjL9vMZ1uumnQeRfoWEu9Hqq5q
LSP4AbBo6vcYx6xUqNPingFS88fDuTjYqQHLIrchFoPD2hW39kv/QAc5JgHPB4iN
GfL/y8BHLLfWPWZyFjrOtxu5gz4X+AvnCLKkMCSWkSTT87vo60/CpvRkKYmdp/pn
iMhqSE6EUQPEqwIcOF6r+BwFThHiN79fwxhdYNdiOjfpnVUIs7M9tOTVD7dZ+y2t
aSuq73zv/DgWmemT/gnUBGdbHGJJL0Ipyb25T2JSZJtFdtblwrt+AuA6fCuDDr20
szOa/h/fH3XyWtJo9ZvcB26cNlmYWDaXGoVZXXzw+Y9q+f7lU1iviEKNxvDB9mKX
GZaAHr5oM3WUlvDa783b3X3yMwLDmkl1mRdCQgdxZ6bfni3yrKlM1BpJN2UGUK39
vm288WUYvIV1QwywKdFOqXDtuqBOTOZ1YaVdRqKydhcNKEk3QhK4SFiuZANO3MB2
iaSTw8hXsf4UrBVsduHB3xI4kt3oSbRv/K6XYudmy0I2iqb6qHr7Z/Z7bcKnJhWm
UkJto4x3mESwPBAtX8gQ0crF3NDaXqdq/MJJiVkurC3x2YPJKFGQRYfOcO6iMRZx
4jiAY3nVgAXnLoaQaB+SZUOoC9+STlUI8fDE9/XZoTzrqSP9m9ukARhmoVSGoaDH
tnIC/qd6xXjT9RKc4DmoLzHtikg220qUmkhsQo+w9LINRTBD7Ra9POtCVl8khJdy
GOtHj0V/CU2HjfJPzs0sjOgoDoXZ8LTPkkzosYoJo1zFMNgeBZsUCSDwa2otQlmd
BplYhnlPlQpqaP/DsjU3JylZJ5ywxg2pYXpLIw8WgP8amne0j35gJGoDro6XVVyj
u77MpmlFboJDErYEs9bnPsNL5ahYOffJTjsfXpoc009sBp3PMd3uS0GxugGIrleo
ok2t/QNQhL+IESHkZdAWv54KKfUMNmTAKYCQpG9YnK/Li75RVmQj7vI36gj3NLz8
44qJP6jkC74A3q2ZJFjJ11nDq8NOCJfyBcUOJHZKCjkShjTo4Y0CvQVOnQMgl8VN
Vm1RpwuPrMN8nw+kHIwMmvzrKzbPz4pTeJQMmQMHhNBIT9hrOMJPhloBXbZFjg5B
kC+EqwjNzOwb6vTbla5FD8H9xE8BTvtQ2NkIux/MMVUGocQ19DnsIFIfmaOIVITG
i4+nqIFsUtXfXMqYs2ULwerp5tEe+tk0BCbIhVIDT5rMKUcyWAOXpjN8eVVXZd0I
bSU0UdsiIgw/asuM+ZV94Ephy73lZw95J3FPFf9vpXrBEXJMOMuTDgUHVBtQ8W0+
5i0+Vgu0krV81M2PGpT+33uJlmivsaVNxUKhQFmKJ/tUo+zXMP9qHp1/eRr7oAiL
9eenL1z9aPk/qluO6k8Ta1DDCThe5kLLHYzFDOJ68tsagjNFvPLvoWNMor6l7P4d
/wxOvFuac82ycaFOGGuVdhcNq4L+wpjtHAtRiEmSY0Gje87g9T3eXOdQ0HOeKrb6
2jZxrqubsz0Egcwf1EJuFlGRcZfiCMHQ5n3kML6d9fuoz5rPSFkipLkoY817sCPi
WGuAg2hvF57Z5UTnbuyzqiZc+NaGO8dRNu6bXZrqnIt7KIcPCEWeDtqmJyj80Jyf
BRnTvZDWnBRTlElscXyFTMRgO43bpblL4nsb5w0OfX0LiRL2eOV6MA78PZsNQCVl
pEbUFsINdwAQMj9zadDCy2nUW9+Nub8hb8rf86vuMZKsZPg7uTQZVP5uM4eJVhrq
lAxmjSHxhPtMUzkt74R+GnA91EpbO6VDgW4Zd/SWmRILGkgisj+cJ+N+8jy0L9DB
MZPUtf+cAXMJ5jhAyHmgrhF2AJkpOaeHHRIcf+Lvd0J72PO9vQIzBdvj7c0HwvWX
Wmw32R/CAwR+ik/KX01R6jOXm+hhWaavUNgqwMM5U0fhQX+Xx0UaPpgM9I1j2Mw5
uLpp9aA/RkwZVE+f1XqQvtl+zeSs/TfmFz3WZSMTfM1WUo7TwcEXTnbpILkYzjQm
FpgKbszqfsXo+Pks+6sD1WYvxNGzj7Wr8dD4x5a3+q24uATunNwr5Crxd8aN234G
3bDOBH84gt+tk8Ec54fHkAs9vL0pc+YKLUkd5wuRaqRtjQA2AFKzVKOtmKOziUZI
XLfK7CDlxdpNfWqEO/EJi+URwvIPNrH6qdBMZsphQnSt/LMq4JLNHteAnr3A1fEM
ahPj55PPTUpTdxK0m6Nq0aUKtMHMLaP72WAi9JmQXDZ+n5iHBOwsqTGnZ8DjzCe0
63GqXbg+0wOs67Gy1lIcwL301lgY+5mm9l9rT0F6vk8twkh1Yjj0FCQIwCcXZDfX
oCfFl5G3Sy7aUVYhcSq0FkkHD4SVlsvpSy49aVoCjHr65SGMpcOK61t8xb0NBAr3
KNSZysnwD4Tpi0ukSsV0h9EiOeGlnsL6AXTitBw/XJc1hf/eb7mna6ytJiWTsoVq
wl6qBXwX65MpP+yh+QMDmi8J2RicNFut0L8FuoRAe2wa2nTPZSYLXkYUaBiHHwJM
V1Pmqoeo/lJ4CJMg7vACvcxycMIET/pYGItu2Ey6ibu+fuZSEgJU3XOkkn45qSxq
7Z11ooXs01RFL+uu0rwRf7Bwc+PDY1zCuViF08ZxgtvYyCYO+LmVgYKk0lwErUxn
4sAbh1iZDXVnDshVqHAVkMWHtXbQCR5EVbLvPR4c/15Ic9FFjpZf7yPDCuFZNChz
zyJCtbKXm1LZDW8AwSzpNpfoQLk9QosSdLdUiznQWSQ1HaCvbJ1AiGYrSKwM6XOx
JOcHX3SGaO8XoCbzbDxQgQeO0gQNgth6kyK5vC/Ra4bsgvocaFNXb3I/H4fbIRsN
OJ0lTNQyKLe3Bt5X81Aff7C6v6ZPbpDCFsaxnAUj/KON97n1fHz+wpIlIIIFtY8A
kGn/6XSCQvjMzYMvRXaRNSSmZ+JmJlfgY29rXBzijjoqXr9uWWWGUOryeB/8/OJG
lcIaCDGveN/EJ7NBpJ2ih/S+BT+HA3Yb6bnkjDDnYg2khTcMdA1NIa3lnWysj4lv
uYKSesJvQQlBv//lzznLyPL0hZ2TaPJ1ClzbuglqFKDpmmzyRU3NvwNH6Cqj0Vd+
vLdZtkizWIgqy7oTTbb4BPU4AaWjhn/spevC7QjsdPkARvZRn4Q1vGzqARgdoyuf
1YvMOGMUsTzbvUb2r/hoRMIRMlsiZda83RDtLA+W2441K6p7aTU/wC2g+cCprJxm
iHKze4cLq+ay7OrgmbZK2l12xk1hCJaaJgw2fZxsqehwE1UBhfLnpPClichoywdw
fNRGddL8CLlASMkFgo2FDnr0BkZ5OlZ4eaKD29g/aH1Ta4pWfCdhIwp30tHmZnUa
hvXF3m/gta8vL53GBK3WFY8CoqNQOSb2MVkoCmKJFyikBmwMjtbcEHNRZbpzwOVR
VSbPEBGlV7T+ToKo3JMwJIbIZpw9nu+xwcFwTjow3QhKCLdHlVrDt0ynF1JtVOrD
CPhMlEAMzBvMeMV/hv58s0KFLfLtJ2Oh7JURp+HsRuGioXOEjiUNrAogPJYPbBGd
YRY+j5/tUepBP1TrQY5/kZ9o8sBVgroFdYR0NVCPLs3p3Ata4Gukt1EEIWGA/t2O
ZEZEYoVa6mgY1WPdd8GXPorp2PSHtK2QE7y5OXgAYlTB5+W2b3V9fsPkmNNX9H8A
pc+e3Z3phhEMMM+SHHMflm9xduY/HwsYMesQuHztGVB7ds+Dj9265tsBh8fxdUX/
ovS+x5T7fzBXk2IQlbeDy7L9na54evDnbSZVK1+bz4+kdtpAeVblGhchhfPtNOIu
Pp9lkqmLF7yE1xOkl0X0qAwZyE5mq61KGzgo1685Lx19/6gzujyfdS++BmaGMHLu
5eZSF1b6wuWwGWNofgT+SF8IubmvEFnnSpKGXcJqFcpigRwMvjZf40twVIUdr8O6
2QIS9AQOp251KkaOfmZeaA4ReFkQA9bRTTKCgIbK4ILw7hUK/sIoWwWZYE/20Lxa
xdNfNs3s9y/WrRkq95rZDa+sziWK8ZMLdSeuwiyXcH2VD+NEmYAg9+asQWQpqD+Y
dfms3Ygh8XGc9t77G3ZtcqAwuWLgBo2BijvSqZqjM4IHiEBOLwmnu8+Kw+DSxAn5
TU8sPj6mu2am3dgBHwbQFW+j6rzn2Em8FrGEcc4besv0xRK7odDjYsZVJpbZLNLE
Ihm9JI9vA6bKHLFYcn7iQMvyNA3y2OK/NkXcL5jRasKuYmcNKML0WnXFUewEObI1
SGDQcYbkynDAJtwPxVRp/b3K9qQIF8qpyJxz6UcNaUVg2BJUB4+PUTHZe3uGuv+U
lJheoezK9Meve6YdYfBD0avaXZ9G9xv9/shqVm3GyfD3pcSbNC6F0EQ7KMx1VNj9
`protect END_PROTECTED
