// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr 25 05:42:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dJKuhuZu8BBLQKWc1nPVYfUH91dDtRiuYbQU28hdEASmxwaVgmGzJrH+x28z8wcC
+dU0QakQyCIlnnR89YGcqLWpLIpxjArSnLU3csYGYT9JCLXGHfFeQpqTfj9bHuRf
oHq5qG9mGB9EJIzorrx2Qg/dHV0huSs8UPzcVsU+XKc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6688)
gg68hJdaV0da4T4tZdz35RdMQP+aRSVXoaMrjVfBTsIc04B69sCt3DVo+JB6Tudm
ueisoVmwIPzsqo81XC2lkRQbNKLj2rJpv3hM+HrDxHSqWpPRoHT0w0tZ0nfJ0x73
P6IxIQev05l5i5ECwuSUC/EStKtYpZiil0IoWtZV1TC/Zb8VuXfGYs/1P0lh+kmi
idB5vpcEq+qRF0tBaGD+UsA6EFoXdniY0miUu/uNW5XwToMIs189MonAU4TDRzcr
3MiPqo2XfUOP4PijZsMrpPnGu8EuKjUm0jyp65iYb9ehhkv5SyA0xjA4a8OEJcFI
QG8MSICUedrM5nQykI+9BavbKxyLigSn15SMrCbDIBO8sddKRPVnmUpzgg308HOr
udAwQzFaBt8GW0DnFSSjf3PnNWiaMp9FV7EpAbVQO8IgAKLPRnntmXjmi0lheJHQ
TjM4W1AA4c9PSYkd4FkoiZ1miCe77V1ttIePAFQvEWxSzcgl3m+I6BlOAl5e4Pq0
BU07aok4pySfxkNIUVqVefAz8oaJhGA/hdz0vhoDiMpLwRn0HEEDiuaVB57Fp93O
/fmfClV/5ReMeHvuG1D/YZ39purQLoJcJzu+a0dvGyOdMx7tlH4H0m7V9ep29E4N
Jo9GqPIjpPjXZfPj4YMBARKXVVKojh2LasHVCmVqk7CocteDvCyLSIE8mj9IrQ31
u+cdLcziPmyxztvYuP4N/pwtvjSL6Al8wRmUEcHc57yXDIHtkNIGXumDHNiY0Pj5
D3Cb0J8m/5RGjHojXKWP1zfa0PRCz53jfhqwvsfvt0wV/06n/uNlPUwjz6G8oZxI
OPRbC0U+OwCl5dRAwLXSBW5uSEc+ITauTc+200uprijC6Tlc3NjWdUhFFYZG+6S+
H6QB5VFH/riP+JVGnxT+nFMCHxgGC05cu3WAIdhd9f7uSeUNxaqFfpPp4wmdj/8t
cB2JzDbMv4/K8To2Dm+3AN1PiEyTw2XyEt4S5oIwFYtcENVWnD+rusFdi+NWxXkA
ECtXR25wT0nRqIPjs6eAr4PIBZjpPGL4nBt9UUDMQo8Dg2Lzz1CbslVpyFic9L0u
rwBjQ5dj//KxyLKw0BJWLAJ2YaQbX7NfHQFR3q4ahw5WK/VCsDFQwN9+SUrs3oKu
cWPStZ89fOzMDv3GozIgLwwD5DAPCu1XEEo9n5St0V6Y5qg0nc93IVCtplYNSVYZ
9wOQl02glxig1LezJwlu70a4uQOhnNFmFpGacxbZ7cISJhJJ/vwu+NlLPkNVreWt
KbP4miX/mdsOtY+th1cdTzc2s7hh8II9hSUO4tIXAXxjhZ1CI9JChuQ+Lp1DmLcw
uHW9Patue0h/1n/OL+cvqAMmnjtN2fp7Cxd8NUgIEZDVihgw+xSJVojyCAk4Oaiv
2NE8OtEloXdOJiUhPWYikH4Dwxls0p5AmrK4j3fnf7nJlthB29mhXtmghfS6LQFJ
EQuIhQ+tSLRaOg8ovhdHDKqszRmKHOg1M/SrePxWc//xstVrVf/L6qlNewSkGaLp
CkJCOfzfvLDPGI77QESiMJVBaF+wm8R96lNkFEmjcN1H1hiCpiaM5m+jh+UEBUwT
EC5SPMIqNFMH1fy4RnSJxO8MOHazltoBceyvfQdQQoQV56962/2xGDFzs4irdGr3
kyRYNpoLrfPmdBzE+KLElghscts0/EU/C6zJYUDTEMn9BHGLCvUZ4o7zy59nNnSs
ulZPMXMblnm8FjwbsJ5vNAS0jpL+dVsZhNcE8jFI4Al4l9FWWObFzvvnx3QgiSYJ
Eu5m4NOXMMlB+5GQj/seId31ZlaxLUEGDra48Yt5agm9tNCABRvXGFJZCnQYshgF
XSgM2vcC3j9gIsstr40rvU3Kl9DNRGyrqsVSWFbLFlMcx3GpHlCebDJlDJGy6/7R
sGpgOqHwTDkzCGJMFyPn/+E4rVQX/Npurp9PNEE+Y2IYLHuRrDzh2AbEByKq9QyV
CLX50yjwQd9LVbokFz7Qaf0ojrfnStwNuzRGymcaCszEVi6rqSTEQBDmHa85FXrI
Iyoe9yQYoVnTViOD+u9ac6GrH8785OD6/t7TJP541zY6DBSJpt+ENVnF6vywJIRg
RMalCO2DPty8FcTFWHUxTggsRn3RxXfTUKmjksGRxi4wFlAQjPcQC2U+7KDBSjmq
DBFuJIhiEHAsD9NsGNrHlETLmcsizPbfIPrRheM6SCwgGTcXKZT+ECdKpOkjEyn4
D0DQe10jgC8JlTDD+A9BU9p4442nM179pyvStccO27o75L3ywkVVOShNATFWLHe1
XKWtaHmkrmroHJMl3Ks9mR8shTI60d9mFfaxASUouui8IYEAG1gj+aCFmrb/pGNR
gnxHWiQvt5ejJXF5GYnOwjNsywNacwURFPXpUJmUt2dQE1dBxLWeL4HQnqDTGKTe
unOv/BzGqEHVAee8pAeFiNkccyeSLL2wiHAMsVzQ7jTpMWRcaMtPkM4v2dhlzP2N
AAfzhdPplSeiO701udZz+/hwux5eotv9yGskQ3E74NdmUDwJv8evP1QHj/apHjDZ
kc5+xwNiLI8Gf5M/yYAYEPGqU/JChLxzBT3dq59GGfNZ3vwrIQi97ybBYPUcpxnP
qqq0WlD4/nVItnSohnSoLmQg1y6ToCFImcYAlbmJmlMIT4l/nE4YZqNgnY6ESswV
f1sMTsh+06qanjZSE8SikwXJLXxs4Y2kbFNW0xGp6d1VSy+gZL16WEXv/HrKO4ob
HLJTBgXeuFXz6xyngRPZ6f34/sS29PIUnocbbs32sYzl+d/5sQZquDzV4w2qP+BD
Es2TawNNONV3ecDB79u/q+FKZLY3niXav2zqqdMzT0tfclgdzVrDMLfILtF2QAvq
nuJvahi6UwR4YmrD67C39+sGgymOWAIhhPzb/Dhw7vAmhaXHPaph0Y2NuLnwspIN
tsKLVJsBwKqw+oRZG0UVCIHDBuCzZhqz577Jc71/GYgrlz8P/dRa02ElifjcNaFj
gxT4r9s5F905KM4CD4aSMhPboNpnzY4IiHNBmZlc6egiBmRUfwLjai8aVKsPznqL
r4NNY9dntBY93C47JR7oXGlJ7sBIcWpITkYfdilPjsUN9hdAtuacG04y0sRml31A
u4OrMGStd6fghzscAMGaxTqNogCRXlHkPyVak+Q9sYmgzy74ioqGDhOfA/gXD90B
2UzJoaaz+ZZ9DpyYx15AW3xgCQoqOg4ykXXcLFNFTTEBb0M+MnY0kJqydZJjDo5S
BRPPseQ92Xl6tYCp+eleA+h3DOLID52dUmPGqkwpvH7qslhiqnrWCGugjO9DXtB6
tX8FHmH5EhaGOXaVnCH8W6CtI14bw+tr6Dys9OB6imCRh21PC4p8vtiLc93CAcpr
VfPXiH9z7ZzME0A8u0dqXX6+1X0M2P2+FeSipSoKsM9JuaLMltlbmktVzlJraNOz
fScxl+GO5sZlnxSGcIgnBV7K54i5TpHn80AYjCG+8MMIZx46xnB0l0lalY2RIRWU
iBQEC7Mb5I5HtO5jGI9BvCnjj8+IucPWoriyfsOGzlzPIiF0NxDkFjiYxSc0rmuN
Acgs46UQXdspGRDKY0gDWw1IiyYKk7WRYEn0BJBGpuRrrQR28irUXOrTHVk1Gxfq
8jXJcpV3Q53BPOytxyjDWvfS3Ro0r056YOqo+2DwJc1tlZFeWQJuVztIMpyL4CjT
r/scGUEFtZutfEyQYbdnhXO9rkJWc+CjdnWDJVE8GwdPX7i4OrWrZ7GhxGoh2CEo
cv5QaiOIEb3UCw2C+bGR2ILSKWNynoPhOuQiGm1kI0AkCYuWfa/IIEuUnFffJGL7
FdLDXTC7BFwDEmhGh4LRxDVM8xkxMj2g3nNPttPcgGzy6PGaaqrucrQ/U8ldNe2F
whe3fX7KHmLY8LZkc5Fx+eBvXQBEjAvJIVPC0nyZtLs/BarZdjwsRG5o+Aa2N0AI
5Rythmp1KspJbp0LuNj30bfRXUurIN3I2e9u+ad/UwCnQhB/Dextlkz93MjpQyff
avp3pVm2ARthk+gNMG5pxcFHEO6hQ6PJGy0CI59ZY+t1I0ny/NddVuhfy3NISSRE
kR8hLz7pYla+WbUPxtiemRbL3ljkv55cdK4383oCq23dUgpf5uoWWQC5PXXfWw7a
S7T28IuBrQU0UR998WiIQ6Hdan7BlNZj2x+Y71XUodXDGzNXU0nYPJVY+NaeVtAy
R2849v9t3MNFYoLSjcsBcVopOWHT9ndIdugqELhmP+5zKBdp1eCfrH5Vjm2pHdsg
JedagfPee+CAv3m37jo0t9icjooxr74ui6wU5DHavcydI6K5q/sIhiaCwSxPgJhj
aIZRkqBaU/mW2PRDE0ZclU7+J+KxUPdC2fAi+wKg4hBTRoKcYAbV5WMvc+J5cMLp
DlS3AmNK6YNV3N0jY3RsSY2ihmgmCfH0iB8Scasp+W/3O0oiFdKKo+I+kZGxJS4m
cIJh/QU2hCbu4Y2+mppmf4XhTiaPpDq50EUbIIu5l4uAEDNgFIR34dw3yxF19QpH
B9cEN2B7aeRjohs3d6l1J3zsUnlyvow5py138zfoOr6cSmPfaI92S+H2Zb3Rsouu
YK5LJXtWXZsJeo2HQcjceglohcloUsx1xcIr6XWv4hF8dMlKuUV//a5wfiz+NwXl
kBrZmd4tgs8KoaZ/rCROA9zs3M1BT5et1ap/w4dKZekycVAxRu0PWeAMhLBOQR9Y
oCaW8JPv+IQfMROVCrYSMvnWTCWKv2w+EN6P9nyuNdBqVsAuBphRin1MfTbS02Nl
NJZiB9jilM4KzX91asNW6UUUKFYQB/Qe0MHJr3kwwPVdD3NzD8c/o8bnHo1P9tgV
1UH4OFKGHRFpRwqwM3IpwPr0eqQoCbNcObNGQT34YlyzvBN8rRp3C1ohaBowyBXX
KJZtKZrmI/+ARtv1xRMIGAIYif78WxRkYwEL0RHYwGr/KXBaeRAIiOQvrqGZGKgG
F1a9KNpbk/eBS4Q7WyKtalDMaCWVGvZQg0iN/g/iS4ZwrqIhgrEpVOCy3/V/hAtz
KnCmaUO4yhlfmsLUdOT8Fq2TNzVCvFoUemyXx4n3eAHvB6ATX5dpUmR2m9JFeCZI
EIigcudQAYP+GB86TvpsIs1/VubeukzwjT9IyG53no5RBqMDR/v7IMRtqpAE6eRK
Ts3hil3JWX0hUodeDRLDDXg6Yk0zgoZEakDN6dg1dCTeBbrMx5EDC2p8VZsrO6qq
EiuOsQ6HoJmk+IyRCdxPEmlohBhSHwikLCDDGdcj9LIMloKcEh/HcP39ilR95OJd
e//myedXrZ9JC14opy6gM8MaSjCEjapTXVxPmAjH8GNOQwRWpyHsCqjK1oNjXRIF
pQuQwGZSEEX5qfSjsC3T/xRd5n+wqzETC3s/EXVebwAvymL+XcLrYlhQ9yOb70NB
ihgrY5FWClVkhiusNzFHHpxz1mxVsFxtlAAOdDS0mdqqV4JFJYwRoKJ5PHQKfgIs
Gv3uAmxMeT+Hep/7M7FuNMom63JU6Obq3PoH1iV6uNAlqP+hPhGjA5adfzaiASgU
WsHcpZhE1Nuhtpj6+lRNqa0DwlXF69P68e1DFXTYza9lbtAiW6TGcMgJvchlMU4D
YN43q79K0uIdekvM7x/+HoyY5mNLBQtBB1mwzbm8wr3pXNcjsQll0TmQOZX3Ukcq
wYIGMHBEUMPnkQobe1n0XpVNM+/AAOxz07Qbt4PHlHwDhMnK4edMkBGUQbEchZOB
llm5DkflkwW9lm5ZPq30PLYror+pItJmm4wCjQQ9P6FQZYDnMh2TWD1OijQW+kQF
AOHYF86gbH57BhyXVESIbwkISm2YEsNn1HDj7NGvzyTrsywL94+dm/B70lIbfr1q
blcp6A51MnBAGPn4Fsy9HmQvPHYL+iqk1QYPp9FPQ4sKz9H7c5RkKdPofzZuTdLP
XmNTkWJF/1bsOb0oIiBzw9Vjph9U+mIAgYtJhMkESDml+gsiEvGd3kNz4KedDXp3
RD35A0wcFbQ/oRsFiasQBuwyJzCLIrjafzaw90tafgHjC07fHEaVvAnIVRcMZpvR
Up0rWRPQgykfK1KCBaLPfs3PTtDz3FNdLhfWE9+esQH1zesoyMesQy1JKyaoaNSR
2UV58QdJf4Afks+aQJ764xH07HIFXnAJp1XbajvCqTudHackmg0Egmg0K1ypMVvH
fabmCRCZt0OaOMobz4GcDjWq2/WWfBD2dZvewNVG0cQ9+B0v1ord2ycdzRU8x1cN
bQ3IVyefLQ6wrJx7GWy4cS6BoELPDI75BbJdS0RuptiNLST5Dt7Ct2AHYSMB2ivS
zDoVqZmS2OCFua76DaPu3aSAX3KYQcNZRGXyfYJxcyTFVTukomtdEJiU2G3IcV0K
5alT1WIO3/gxNFSk0uysNVM+BNSqrPRKtb2UVy545WtPZjSbEVtO6DEFIbwxxDcX
WCus35+4CxhWteVGNqSfkz8QAzQVBg8KfB9e3gproWTdN2mRFFHXHwlyfttM6WT6
KOoiUhSGPWTtEZgZDztkjdg+B/J3R3dTFxY/gs827JGPFhlKrlUUG3WDBdJiiIz3
wLCw/ktlaZq/0Y9rKRFCOX7Ntmfq54HmPiJCk929s9HIoPxcoca/D+aJny1Gdl/j
G/p2/5U1wY77qSHpIsWdct+J/56j22orohgPNIRH7kh51Ulvoy4SJOv1bnf8aHVh
/yDh1dmOyZSnliF7rSvfGCA+j81mtDwHXc4B/YxlCegX01HQrBSA01x2WVWonZQS
Z8FNLHOpnX+f8lVzCFcUvp/PgF9lvhpmJ9LKukmx4deEYGUyFYMJoMgCpfHOm5nA
/KlKIB59xzd/1uxd90+Ezhj88Rk/+691EmhuU3u4j1axmBB/HhrPzc6m7Ntw97If
8DmypzHOrF8hS8qe7CU20cHXwKPR0zkB/vsR1Ql05a1M1Y7j15Ltd7jJVv2Bb+XJ
DBgPH65hL1pCNIn/wHJvtVs/qHcoVTq5AK264IJyeuQQ6cwxRzET64SDR4nTzKAw
Vn+731mQ3uV9vt/pOAWgRIDR2KnKHEhcBVqKfdSO4BkhbHDWJKVJ6/pOJzfgzTIJ
3jJMzw8aW7d9tQkbx4HSditu/s7+Dgc6ENC6pWybpGM9h1zgTAgX4Ozkf5Ko3WkR
aGJt6LwiCXObd/OIPFQXPVhbxh4CHrGhkbQx+u+w93jqHGVckeFu50vQcYjNVJHt
KnDI3ljmYC8JeXtjoK4Ck3zU6l/OMDaZSSQzoYTid0TWV6A9lAEeoXaeC6PwaVJx
fXkvDvH0hP3y31M4vG88whsAej5e6mgMk0ypRfY7GG1mShE7O/byElFR56o+UUAJ
FO8OTRBLg+7Rpawu4nwxHlsto6EEkfQIw7/DAFhkxuNRWywYG0XXOyGqErC+qPWW
9o7mjwSwtD2WIgpZkoaLoT8HlOodkXm75xejJ1GJ06lBwfhN//+pwx9C4olIJUzW
H2RcxxNe7QGcIqzy2bwXPZ6eUdzCQXEJnkE0qc4NbJL+yOsB9SWEf5EzLZqrzXfR
aQFWHjWmz1cEUbty9cI1G2222Ka8gNvAM90+ierI0+HlpB+2T04vyEdzh9fD/A/c
E0poj37cnypv+mh+pXjXSP3Q4S4KJBLYw0dHa+mhTEKoqWsPDqhBkZC6u51HwjUW
NhFGSqbHOYJPzNFWOfVCvYtyOlsiNi0W2r810JLhuXp+M22jjNYIvWYOkJrs1QcI
8lVBSLHo9aLr7+N4nOVR1K+lLvdm3YGL1WypKTz20EpTv0NlL45B8ldIpCRaWqun
gEqhi74Y13w72ivN9u28jyAkfP+BTyrtQ3saG0L5QmmDVxFtuvSzuW/RodJXo9zP
10FFMX1rY7A3RKlX2kF93OkeaKDgv86t3P7+qN3+y7ZWf/FP15zBn5wq6JtdDNrt
uZ+GP5WlxqckeTLi26q+6po04oRDNj2SSPAPiszfML+6sbfxIHFdopLj1XxYat+e
njB6k9cJPS5KyvfSd+ffzZoJIQAtwws1a9kQM9dWPwuxQMmtqnjBTMSsSTPTigrl
CUtmHkK3k9n9RqaQP1GJ/rcBh3C4Ke1cPU5Ct/BvnfWdpnkhz+2eIJTd7IieiibN
D1SRuqmTyhYjsYVlXA0TG1MujfGOJ7xpyigUVFIpBj3ap46ynZaNDluP5aJqFxqq
Ok2tyMgNiiRVF8Wke9+subsKbvl3kYRIlWyQjQ4i0wKko8mn5ZhdG1G0rIgPC00y
gnDco1+DW9UJHiyIPVb3ODIipLVJQHBPTf6VkiQUAFUa13u6B8fwbGBpemdv54Ee
Bp2OEYqBK2DPsdNBZ8gAcixXgWExJoMIzGYCXUTj2C2Zo40aGuH66ho1jBbDfVoQ
aVcmpbrjud9KaaoAQxAr9SrGcqSFRMB6ySYTSbCT0MWhr7pdwA26K+9VaWfIHaXS
TGW16FXlLk/3Xts/tORY0GdI3KiWYo+7siBgqs9b2nqt9zMcnIYOTYl9ABUTRc9b
nqSjh3a4kK8Al3kMGoZXxcKf0WcoCnC0R+yykNi5Ee5FjW9kLZg8HWVjUn3WOXQY
ulhwLCoxtbxILdKzIt+JssMwcKyLFMl+wVV3hUq1YzxCQJjvdMFOeSfkKX+ls/9I
U/V4bZG377WlA7Z91cUBEGA6cTeM++f8AnucDLIWwgVBw5WAmvSmRXOdc3jxBC8R
YOU18nSLhQ4cgpcSY1yagWXqPKVkmx1c+4FJQw8eESatqlSc5QJceNNuWStwuuGA
AEq0Wjx0FUD7D0zAoBvfx9wJEoB8fqTn/ZK5zGGh55f/S1zLUA7WDzGPlFF1f7Gb
S5S/V+KW/OqG6A1EkshzFRgGsGnixm0MEIF+CHHRc0GlvJAvlrc3bVc8F/ZWtY76
G22B2YG7T0iqYz3/r0jOUQ==
`pragma protect end_protected
