`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tGSd/1Kdec5p3Yd6rfHoOYdQj1j5tEgP9KEU8+kguPSWVZkbEEWy3cHdlWTDsE2I
VDVHqmRW+wadTilcMKaq8bcNkyholdg0Ho3WswKe0Pf3B54bxJzloS8QE2PYmRUt
9Ks8LhZE6dLmEDi0jZ5WmpbdfStmjxMysVpcAEmXAnUO8aXNG8VRRo8Rp1GG/7Yc
k61UvPPfNt+rp3LTB1lot1RUVmvxtuKjbrmVJwsfyEqvcBA8tBPW5w+oh+h3cjXq
2Zfbu+DbapWCKOoeXmVU+0Zp11aD0wNih0HUR78WxnEEpQv5nrk9DImj2GZhfzTf
n5dy2iEZnXoRwqRQCYs8lUDclOnm0RlvijBA/elMLNut/K+U2KkW5lPHHQ6l4MQU
+YJnSDDnXfq3juKgw8QSTojuMr4KOKMbhs4Ktd6A6KlkUENNNlQQ8DV9RZGg6Lmw
GkhOBacF6CuGHBjTLDeTFTHo/n96LwIOfQ+kOSQyGwcOyM3KEjPeiv711PD6f9mq
zveb7m26yG67mg1eH5h71zENhzRSHmZ+dze1ysIuOqKf6RFvJx9fprXvmRHI3ooQ
5xq4LGQK7SfcJqTiQo9ubm5VzgSuH0bXbyb2Oo02Q7TvNsX9+D855gzZsn/fvCIy
6lYWazBhEuiNhXYXvG+9rdKLJvJhNQU+R5Hoo9Q2JlAIAvWHK+HK/GP7O/MxqKee
bMHqCWHs+Rsa0jNylUMhogL8sziffvsB5ufjSqDdZBb++tOYOGkMzixuPJ287Nqa
119SVBk5Ft7PRIo/Yrf9PQT9bop7tvkrgdd2/tr+e6BA0Au0GchTn4QVF8eqG/GR
sCl3BtdzH7InZoIXSBMniCZguMyrXI5tp5m6+TkJmkUc2yy5ZYACfPsM8L/Huhiw
/QkcCQHq9wQf7CAd4L0GuLvbmKuboL0y9tFhsO1814tbC60B783KysFv/rYVbJ99
fLSSrrpfSDtWSiVDKUtZJVjUpnL0+tUahH65rHyCFHfDoox6O2UjLGZ4J/ZPFTtu
tzE1wQf4m+kCzg34eOKmQfxn+XSqW0ylq79MfMTl4m0crwE+BTmLMrjzyomuv2pY
8OkXNrRVJcs4wFR3kJpeieh76hl7HoeLYVzQ9wHGgC1SvEJtmW0S25rQhwlu2B3j
vtY9LqSjCbmeZQHcGBgSKJRk7NyEPodEKg1roZS5zKlAVTby+6hC3+1Tob9zznxK
DVfQ3X0V8sj9Udmhq4oqfNbee2nGICSCCKAdO3L6BOpSOAGOx/KJbAjmfNxBrWlr
OBkOat6ZNRCdpwCNLZz4voa0VJ3aEBvxFk6evk0xgeTR/U84nxOApFbPaBL98ALx
qruXSgUAy8gQ/Xh5Al3Wltg6cSwlrwWs0aFK5v8nwHEaRV5QFL852EkB1Ei8jGxU
bRWj57/9joCS+N1eburrUQVdkDJPzMJTtg/YUui99szZtjbquuo0X4cGD9n+gJal
5SHl1TI548aWCUHoj6t9W4X5ktrrgCSFSHrjub+BDJ50VsgHsoLAQv+JxgRC7gX2
7I9EF7ULTvCFVKB8LuI3ZEomlHJrbR/PE35a61V2dn9rHjikihECD54715mB/VNC
so4SZcBEdbATAQzHBF5+qNdpGZ1uIiRm9ZwdZbX0THWczHqDWyGknCvsKsAz6FK6
HrBLXKEbvCzQ8hg//TV1tpRYblIST3B9BH72MUmdTf4FMwu97UxJbeJSyKquVGOO
Ot7zcFMFEH260an4nQ8RO9oi+5iI5BXNQ4IGkaUkh8ZMqFHwvme1KORC8gZfDWIw
2C1vhkQ44cbCU1i4ZrCNGlHZkoDD5qTIOnSaXhpv/bIPkgT3ttfacQ+Ug8gO6/JV
o1rgMR7qK7lm12RsM2BG6BDONtlFHAIF7lHQliAkzk4ApD+9Lj+EW3kbGHA6WIOR
aAI26cWHbhLwEq4BlTYJw39jUptXBTkFv64EdfvzxtmyBF8pnYsgq1gQPzJqNVQY
6EHoqm0Kc/m53xvsc7X+5n/JS8iUCKh4+lfNo3WqXGW7t8qutyQHIaLuXWbyr9Ya
znlQhQY8UCm7j/NXRVcyAWQ4HCKZ9zMsZQgfMsDggOMp0nQF1Rxd2GsDSKoZOAFg
cLaOR8Dq5wwwLQOcGxOC/kBkGlePt7cXBPCp+I80TeSjYflI97BAAqV68Wv6yzFk
D4Dvk/AF1bePn5/BAbIzbiakhJQt2jN6FMeNMXYtctSvibdLHAX7kSgG3yFH7Wei
d3Er8x5MKVF3olWnAt3oHxaNymJ1VlkOgd3UME09fjVf+uxEKsTJu9vjoknAC3o5
lp3cZ3zqmKtHwhgUnoBl5FaonEB6Dv0lno2VPy1JBEjekwJn2oNgBAGWB54Kor1L
JHPFwlVfdvzpuYNI4XhB5ujGA/J7JrmMyxAdK9mnd8ItfDL2eI9GFV1owf6CQSOy
7jKVC1KZ/E5Kt5PHjUmf8k6tsI8c/3Ty6cV/IO/Zh0kwIx7xiU+x0oQo3QQ71NbE
mZGvmD0SFoPdyBXhu6DCCb2L32llzmD0JHclPQtKE8SEsVZ1UN7kUl76YWUGVkrq
Y4pq364+zGUy7N7ul7sFDwLN9xa6+eezTRhc4hFfngBf5nPQBFavpDHebdmHjN9y
f7a6s2cd5dXhHds/TgKswJFAmAgvilJO4UEi5+tcnE+8yjw7oXO+IrqUdBok62HG
1X47Mk7Qox4OfnRD3Hqcy5wtAzhp2+/fKbTsEixBD7asdXjV7kdtBrcKJMKRTwxc
1DlZVAxBWBamBh/IA0SAMOSmBccVFgdp2fZGRBVDdwx8QSvc+bbxSp/8ovctb8nN
fBRuBiA3FWoUuckNXAnsaRdK1qg4gY4uHXaZdwhtkLlmKPogMJ+HKxtE5jAnvBQm
gatYZkHuDa5z7b3EmqpLv88CV3StahQzKiLwvrnNqmks2Bc+0S+ia23ochczPMFT
JxWWscgVQ0fdsKcGzYhJccvY+xMuaoHrmB0/HzedxBpKe9B6PwxOwAlxAPV7h/+J
/aAxnqjRiSvRhKercFkeZ90qefL7nfGHyWrmBT5hHayUy/H7rPmq47BbFIflDkup
gkjEpxZDQk6nvE74YncosZqadpwm7Fw9dXW6rkPfRT/ro7nWdR+ITrsRP5x8tmuU
JD2F62wRDn6BpaAXDEfvYkFj8UQKBrPSIa0gpzhF+NS+agMEw+CV8uV7MmBAcqot
953QWWFSlnX9sbrTdweuovZEVB04jo720hk7/srkgLV2VGIJJOlhQUru/Zq1iP0/
Q0pYKgUCKZ3xyvfW+UqLVu/4SLQcislDIHuYxL8A/1nTB6hzsxeBMGesS/nkQo38
aPKRyPMG8uA9vI7wVl8hmQj0KbuRz6n+CXl2JJqmYqb3squB3VfOr7q/yoUnPs5P
ianZDijvEM9GHE0E/VcltlPlaO3el0YlvvXF7eSQ/q3zQaYWrSzLPGYmnmOww8fD
W5UFgZfY51yli/l1SgkkdQvPU8R2v0CxiOagh64ZyqZBvQu/JfPg3WSXqFY3Sxpv
KD8JoM55G0xDIe2XU03wj0RqI0Rr21y4JvSUoC40PSvFr1SXoYHGudm3ZzGt0hVa
gGMMiWqBbOsCTjY7Y08q2IpyuR1WS/LgJCm7k6+7CSJHQgBLfDWlHB37WB0RAqCZ
32i6osPrGearTcQtztnPd2a6Bl4HQHZea7riyKa6Um5vNnxrax9lLG76mk6jVoGA
inVWQ7k6JBCWfRD2m8AuItkxe3kcHSjPUPOQPqJ9u9zbGFvjuAeILIt7VR5LyR0M
YgHr//IPY+FnDBnJ+qmdO2bRlk5a6vwqBkwOMbIlG8j873qGIahGhiOF4rIIZl9o
WbCXDrbzT1c4s8L4F6HnePqtuKnjAEYwoLhAZ62420tZfxcaBijRBM2R3u5G7l+P
0oIF5lPwgj2k/lzFvo1iXtXfZ89l2KU/U32EH8PrX33KKTCW0KREljxBHDq3oS70
65KYVUPmQZX6V9j9qyXWBSIO0r+7pyHLRHrB4/WHBzfiGEokUvEoQ9eBcl8rTVHo
VSVw9R+yBIvfsosLDD/is2gcdyz3hD1555dgc59vWYjNfBCRxDDJlDZEy3NQPZiD
+fLyB97ZBCwGtyHkWTA9xuo6tfH7m1i5UjWh1J8CYImuqxaILUQ10wepKaQvVM7V
MXeJGxyGN6OeHoneSqNgu3IZ624Vquh5oIvC0ziD+SOxA3lRDPHtSvZMxtwTykM4
mdBVIHbY+CAxgVkq8Y6TgHxzTNjVTjEyrUok1PLYgcH16s8yoQprILp4W4vwGLM+
2YnpgB9/mvBwGlH5U4YH5GfsQ1ih4tWhsx2M4yequy14T741gj5rP0JcrJxemkZ3
U/QRuQcT5PYr4jMdEBOG0bz4odE3egqRGboByvL34T5P45gRvU3DlpRgboDP9fRz
H1FfzXXu2Bhq06j+gmCSK8CJ7iW9BZF1VYllJk68pMtsE/+Ojdf5waJk9mi5bFcS
RSfPUXYjJ/IKbzwsvKishiOeLZhVLMiLjOmGi/eqLppeEUmn92G6+L/VkL6Cl1Ra
oDsHRCzIFGIha6PbIQbMXoG2TskiqrqGFUQ2KcaxEtFsHuZe0JWeLffdWx7/7D4y
dGMZOaiXTTqKI+OFJYpb00jrkGb9HOSqhW6cw/xDIMeJzNIpBQrAeDiEgiLUMfim
9uaPRNg4/Wf5hh8am/ytLCXl0kJwYzPMV2zZmx+wdw4RZx79DQMwXaBtcBV9Z2VQ
rPSBDiMzwC+oWRkixstK50/UrvutSVouosi7vnPnBHS9IsFPiPWcrcP1mMICZsOT
GQsdB4uQy2SoKzrZqMrDrM0/y83WPWDuz+4k68osiI63c/8wazUJUuhjai5XWvvE
NUZh/FruHSLndfOEBwDwCZM11cR4HiQcy/HJIQiqlK9SjUBq4E60JkQgU/3O514x
heNr4JQM3G3pNrCLa/hCUc7mmzc6OV+zjsXvKug4gp4icgM3bg8SaTUJycrUbeYZ
1BvuHwDUhJxOZYXiEAti+hSbQQjP5wxKkcWXu0Zl4FPeAhFi+i7Z+o+8P33K+eKp
lKJgvDaB3cSzAmNhLGDFtrGqtLsVx8/65B466TQm7C4Oqhs3e536e901IYWsGamr
oCgJI5wBYEoneeZv1Tb99p10ls9yea5iKQPdD8djvWv8uKAaE9O5svDxh3m6DllF
NgfOBrerKNEfnP0WajWysVLJG8sEq/Kqzel4E4XNTKCB68qCE8sJitQbJdIpVnY3
OM/CqOUP/100rFMwJfZ7gvUkiBXo6wMdXpU7A29tKFSJqC1fV7TnVWNhgUQWyODl
4HlEeYT5KMmu4uPTjX6Vlk0+lBOIImzciU2sVfMZpntuLH7HYklcHLhdbGIpUu/b
Ahb1JMUjkY2kRb4ATHfrc6vzB7CaUBSmjNvb0EpD1zBgtomrVPDhJ9RuaXtD0YVJ
Th81k4+xLKP8PUMdQdLTh9mq3RH1EXM3qmJp8NyjESTULU+usQEYgoN9FPELn/5+
uv9ZhhoZFQZ3RAPqockLr06rtRt4o9xYZFjpHWlYut0IyyISYUYgVGGqzvxVZBcE
zKx1BjZlvXWbTATH3GSA/N4osrXAs9ApOhlVXtId0AnGUlYOOYXYJxOUzDJ4IWt7
0MBmGYlbuAM2QZ+JfDosQezHRaiP+NQCiDcunjCAMohh4YeshNC+Rd1DtlpbhLrS
zIognU4mBtnUMB2Vs2sDujl3Az3iFGAXMbF6PafLZrZ7fL64KvRp50fkUo5nNX6J
WjCHWkM3dpyOjgeKQZKSuvzZPXtmp/pumezOApAjV5ZYhuWYMSlR1xMcA3UzLtts
Te801NOZJLsQVmbpBWDcfyfcXGQ7wBaG59wdZsTCUoOvkpGXu25eNZKrMdvkjL9r
32iGSF52zpU5ISB1v6+Ark4S8mPDbd2exgTWPB5r5rI5Ia0KJ7UT79oUI+YIWggX
bEX62lwtD05WXjcdyGN8tBSm5Sewe+iSohnfLN5+FZEqWAri31WwWbKAW5OZqEDF
Jg8kqV3dd8oaiVxsoG7iWNfGL+cD2Adoln26cBrR/u5U2DpHOs+cwIZKmuy/3ksK
Wiu8gQB8G/rzFxt6AJiq2QcVvLVlJW9FMvd+DSFNtakAOMVcvBFO3T8mCMhUya0K
DLkK2ocR4cnf7epJF6KaPsEEAcmSKKJ99pD4ldBZqBZIoyAh7i/7K5A/zXyM444s
k1wfd0/7M6DMwKNAGH3U++LU6Kw9Ol4owQk2L0AbXF2WHS7zhg94Y9of8raoJGK9
sz92MeWLDKXb7VQATLhE/pIqQemCqQxxAhchDqpwzh3NLjOfmNFYQjAlTr3SAUFA
bFauQJ5Go8ELoZEzQnVxdhg/ZzhUgz3ctAkFDD4h6khfOuNoRF3DauFsE1wDfDGN
9WEndSClsE2W7sderirtwfyNWH5gWRWXCkqEpSlz/7tWikp7JB96oA/2irxrslyP
1N5foKjyE7MAYyzE53m8QQ1ROXYX4+WtM83teYQVIlPTER6easl5OqYJTsaBqTAx
IQbilqI/uZy6GgbHTlsg5E19jYmE+C2/ZbOiNT/0OYj2V/O8/H1J657o7/X8/uuR
Ss4VgyM284VOebhfQdqgpcTzABbNbkW8Xi0hjBafsGmQdXkjXiGIJU/279XwCJfY
H4iS9LqmN6nLksImW7NFrlEyURpvgSpXuYGHfO0bu4frPtxBZx9UFGFpf+Cb1haV
70mOBVs+bRuWpRwER3pmYauyxA2LpQr6DpUHL0UY6UzEKXbgztWPtU3us2RgS6FP
pztRbTJDpxieRcHIvrIwyKxTqklc6NbS8EoqF1ggM2GIkUUhVSLGVtUuTAAnM3Lu
GQEjZv5NSyJk0zOhslSptQy7rqSangbF18mXhuiVMjG71DdkZjQlm6eEWQ2xjxRy
wAd1wKjamZAtZChDiBtlE0V2QDOxZWJJO3c20gckmbpnlOY85QU9sS8dDxM59FP9
1bk3BZ2zsg/gEclawdyJdp37qv6jI1FFWCcru50ZLuYFrbAqQ470M+8ae+nNd6qA
IRZpUdRNa8oYqp3g2P5a9fu8hjVRZeP/jxNg7+8CpGG6CBHlGI5bgPNaeiUUnBIH
42UKbG/Mj8gI7w6OoMlyNpeFoZQxurbu6hrb2cxuzBTgC/ZrlPrmI2SkA6YMM0FD
C3OT2k5iwu7j8KOggJkJ5LKQyu1QZOQMcZllkpcWbg8s7zb/k7eCryJZx4GshyGc
a/R1DQlbI3TSKg1fIy9diZxOzYrf7WTOAHK3s1syPfbTbwMRzQEObGdA4OSc6JXs
cK0b3+pMHHSA+nOumrQNmmShlSukGRaKSBWDGK2sQGKE/v/QCiw9anHz8OJUsTnf
ezJs3zRBqhRejOZ58YURlkLKBClyRSlJbsooSpWS3yvZxhgF4rZ8gLBSGfBqLMfW
B77dU9IUKROGYaFu2zUbFSNnkSnPzn5Ym58iohrq09UbKHl6s2hI3R07TZhIFSrq
p4MXoc8Ynd7u15d994jLUGbOBRwThGFrM4X04jeUalk4cVH0LmCYCbUy3RMF/ee5
PqlipRCS5eCl/R4n+1UX1Xu+5kxrPfSdKZ4njJyEMnRYc9cmN6XnOv0q+OblZVef
cyObipQ3os/lwESVD1uuOcq9EORv/u42AO6TOGluKmEMG+u7xLkTKhte59DsaD6L
USFN4D4+OHXeo4IU4DttGq9BmtddBgHpua532wZNlAqrU02RJuPcS93stNWS5y1p
Oy+EwnF/1vcBLCnSe0tZTOdy4VwmFY9/RcTRhwc54e+CgAiCa4LiX7vkAOmuryFn
roYRwvQo2wlWy+PZR3YZrmPA0QkGzsKZ8eDBiGe/k+HsVzBftMklFY6oDLKhol8p
ZHKkIoUvJoyA5mKkpSQgHv80uARI5HAf/sk0x093C4KbdToVtNAmmltj85moEmpM
YDgph4QMWTBFqdAhC0Cik6xGRc9LwpqTXkrfjjQl0CgVnzNrfD4uKjqiF+5A0YiZ
vozpM6jR/XnqIsJ0pnnEzVd+zjygBG/R79MO7PNhMUtTQ4MjNO0zLRoKb3k4jnw+
Fa6JazhsnCMKZ259eVJQF094qH6lLLDN1vJFvoJAne9r8JKO3cRLNzc2Yr4Ryo7H
+KC1N1SUFzg3U5ztyNZ/i6+ZAPtgXeUEPEnEl2jga0pqLnUiM2X0NXMDXrdPZzY8
XA+c1rZmFNAVGLCLUBaJ53qRgzjO3IGSfzOcwKobxSOOfGujZQCe+GHuj41DIU6A
xYnfZ8Rzi45BZf4Wirssvr6goL5+8Q+CDd6K4VaAIcuZozC8++QBCihqz54UbpPs
xkMndtRqfFzxUKUcc/WQG97/+sCgAx9Kg19MpMHRozdE1rVY/P7X9Q3015Agdin9
6OEdtX7X3Ucf/SxTPePRPYZQHhYag/tlSjs5oiJyrro/to1eQil6U4uZMdres2Us
mkz+bH6HC4L3wlwd6JDH3Ng45VWit1076WRCKH3MNfTro7YLIobm8XN3MRmyA3T3
UwaWVUiAoopY9g8Y4qssNbwI4Z/p0ZK2HeZ+vmjW4LZ1aMNQMgBHVc1dcJW/s872
5M3OqzVr5dYVO+TFi5G7mO3eY2pIOZxiJ5LtMK7E7bO48HVw/R70CpbT2P9zVlCI
jsKjeyaUvQBnku8hLuPpNFsFXwoXzrGTLwl/HFDrNMx3/zyFkZ4+oQC5PyNr9eCH
kZ1ebZ99+/bPyCHzG5i+gsDg2dnVSqqDQ2FE/+PTtx78lAkOTY6zLiwu8XtC856W
l6jvbGd3M2fZM1k6NP/Zn6H9cX1GnRWCWXdRGKHxbrg00DuMJf5Kgp3N6zvWLsmT
wpp6WQ1g+ObYqHM0t4qoBfStRx0h89fl9QtFYpMw7jojII52Ok+Naifa3DoaaIKZ
YUGaFoJX6ZzTPst0FxLpjd5M+iV4PxxMSzDkxxV1nytlzF/JD/OQtDmbisLkXlIc
cssWTvkpnRFc7s5NzpIdQLHdIPmBzFXOWQU7MGQ+6/8q0ZCIS793OQZ5ZlGx70Kh
s4IigN6cSZGrzSsr4mKArZdugDebesTaBT1JxdEv52vanrzLfQxlYI4dfW/teuBV
eQ0c02jRwPpLx1CNFBe+i1W47ZHvtmzBppxOcUX1Lgzy/0BEQbS4i0P+MG4fxCag
AGW9gn8oF4sk2aktZGvp/HCUrHumDAenBpHE52AjCIBMxFFhQbrB/P3xmG27e8Zg
PwIqi58MicXiiZOdwvC0yW+rjfhbqS7b+2sE7EQbqQpexSnsSKQE9+g0pd9mEA5t
FEgpp1ZcEbiWndGXnXgnLpC3JJrUSeKr/o/f90uugAhvSkPO5cIWtGO/oh3k3785
xEOjrU5jelOCOGe+yZiIwL5JeiKATHMNdLouzQU+ZY3iU8TX4m4dWSVI2tYbGSCR
KZO9GcPRSmAq/FvFreXtoAqLiACSdHcLMlmPhJnGlwVV2XKXV3wMqlDInPdj38oS
r1RfwMBWQskfWoMEYZaeAAhF8DNhyfFIViWhSlbQ8ahN9BWm+7550wKagrJqtQPG
nn0jwHQYdvLKz2ZKkwgE06wor2z4D13hSKVoOoTpWpWOjNTrljisrDU1GbnNRlWZ
TJ+j7yAdHqd3UqtOifIADVKYtbFOTjFD8E4amKghLU8byGHIFYg4ja9g6fMuo1a2
Yvi86/G13zyWAWkeTBuAH0mI1tZxhRdW5hx2nZ5QBzW8KpUrCNSy5XkzO+/hLlxq
y2teKLkPEpdI0hctG1Bu+yJgmeKwBVejXS64sZ6LlumDsLwQjLdjBqcEEiXx8+Ad
hT/SaeVuWvF32nXzl4gQMc01h4twpHDavuurkxYg0d1sH1qspxPPI6srLU6j/VSo
AUk5RohLZWOC+Bbc0L55m4/SfF4Qv7aLhzHwBV+mYEVpBHSFmGg+oJbevi0mXeYV
W1f2mqjsRLjemR6Dx7uHRhYj8Qag29vtYU5ruNurPqjiV6eFb3EzMR9ZuCPSUVQk
qwyWtjzLOKreCBRHh8oGGXgosAnKdFPMMvebXLS3nJnXqsStWDXajEcDgA7/Pje2
Mjoux6RT3Y6BUa2T5Ln9GFmhRrhIEESxcH+/P8zVAYWn7dCF0LqZ+BhFUYA7455M
t+B3ffSS8G4ZTgl3s944hlY8YlGKeIUDWJB3JZYIyOOavH8MFz1oCo3ByrdaYoio
2ijCxrkS9dx2oNrYDqB4DDOyvXMWuUKMptkBGL57eftzvT0tuLUCtO8E1oLJD0SY
zpRRmi/VvwBF/tnHScw2T+YMqPqKJnN5Y1UkA8w9tpJuxVuqCVE7Mn1OdwYrUQp+
PlqMCpfodl9YcmW+ioe25bFY3b2Aur058MHmuhBDUFhzIoVu0CpblfpIBj45fx2R
0Eu8GXm/Tn5/BQQrn2gvURdCBl6TyXybm+M9J9f64HDWT8O84hTOwSWtd4Q8DnMd
2oQnButWCd8KL4/rtNPezoXLTcvWCvWo31ZPNQL4yDtcbnhdDsU05jiTG61akkXW
HR7KmTN3Rc9blWylnq4stymvFo8t/C92wM1z8YeX/TpZR+OUAvlmc9LNdzz6Wt8X
+Iwtkt7hoY65KsQ7i+ptbIDQ14Nod8DHCmcXddTivrnHn5p59ZddUuQyxHcHsXeZ
DGgTvLs7Kp0imdob8BOP/BnffVQFXMvHd4Nt2ZGaczVDNAtP9PaOen5nl5JoS0A5
KwOx3xPYc8Hd3UZdqJDS/rqxhwNttta9tZ1G+L4VeTbmKxKcgf+eFq6ngzOzzioE
UARtWpfotS6NXG7g4mMChX8eU7fnyWVce36BYkL+L9wwQ466eRGVCa9xORNCT1pu
shSRXBdgAhEZBGu3CzW/UcBHfHQ5TMis08jNFClDqnmVRqu4GoiCTRkbCM4qYQpR
hBQlxqZEpMNzXXQvQlMZVwUiiHRaftbJh02KLGJu/RVDVxE/hXVlchEy0mVUJNkV
dcBrVtUZjMVQG/gcoieGMDam6+qkqSWPGsTwRlkrnwFkNt4hjQ0al8T8KUFiqHWR
5R+y2NGnLhwBxyXntyZl3xPj2DRKiQzibxYgXnHPMB5VlypzYm/T9SpC7PETJZce
7Kfq981XQu0I28ED4g6ITHPYrHMhHSbuqSXZp13t7n1PMBucYvJdZ67yCnK7yBXZ
TQlCwF481jy7cnODLSGI4anCgMzd4RmYlUf85qv4LuTauOOFEiYcbEyzrL4MnldY
C25c9X7TCdpo/lhjCXCUgmnSqsDbcRyOtRXzoIaNVr+OWB7i/2Uv3zj2JpUx125M
VELYxwSgo/241QzJNVqcRres9vnf0QRDOkhhsnCAbWYjWlUDpGTxcdda1NmgfCkA
N7ah6Uh6c73S+6z4jdXmVI4C3xHgBQl+nxvaUaiJbc8rYTIZjljZVU2jTsJIIg0i
12mzl275xh+wTaN0wjE9i1Ati0YwnX2GPOCj2BD9e8s4AzRvZiCRmj0A3mBdnRrN
cex63dbg3MBJtWYOeAK+eYoILZ70s5QxwfvNhbH0mdMxkNPp6htxY5Xt7Ho57C5h
n60uxTMv1IXm3w6casDx7grxI7rw5R4akhLMydzXUW27sGe/yTU7NdWkWJvP/FJq
LNQ4/azxX6Nk3AEbzjPgUWu+sW+7oCA7vSoQQGPdVu/hgZ8pKAPQibHtgk3dvwCM
cMT5fZa+fKscSKco7x238Qe7H8dzTr7gK2UHTEKmOKilx/27duNpWiVu+B8RT+ri
YfHCgJMe2s7rHl2GP6/x8IP/v0VcysAY8o1rpt9fDzWVH3O9tOQqlTqZynvR5oLc
5HoSiyVB5DD4rzNtGn2R/Nt+CsDhWspm02jCyUAINoXJYPWFV/x1eP51G++BpduM
Eye6liIMsTSbe/YT6WD4KB/LUu6wqTwRwyOp72InTijLxBf/g69cRyh9xpp59f1F
ap4G+wwdsfqONxXWDxm8Dh067qd3Xcy3O2U9qjX0mBmUKvq5Un9BnOkLP8VNstA7
u/HbPBRVrKll5ivwvt8dH5s3SFudbfVQ6pIB1QoN1I5dDNeBRH3TYivHDnm9uHoY
gN+70srEk4zh06UeKUDQWEJlzJRH3yUfHb+dXgClsOu0Nwf8tl7Rst7akxKXMBct
38kKfvXgvzhNFEjtUCBLMy+N9suzlPVszboo6e/lrZ+4T+cYN1st4FtxPfatLcFA
tUixZNi4ovdYedxy1jpM8Efr+KxoPoKWIASdo1Hfwki5zqLFqRsRRG2+rSYRAb9y
xPqAZNvGnGtPK8WFHuSSgVtble+5KQKVxQ7KuXwuk/I=
`protect END_PROTECTED
