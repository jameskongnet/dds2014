`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y06dCXcoUb61fJ8QONwBJgeX2YLJfzs2O+X/yOcs6mY7t+qgdw5XATEDGzK6LXRQ
RHOggzt4jbJuBpqCoC2eiZYvZoTaYoXUZcxMlX56mJ+gOTP/2PHTCV6OTRnGxQaF
ORba8w2/zn45L6dM52HtMINFFFvja1zFw5Gdrrt0caQuvzLtdzpo4Pj7G6ZKHpst
rg9WnfCpC6bDlkuaGmL8mMyQ/mkZxd01nanByGAIpH3HAEbf3HCI+iQLMM6M7WOB
onGLUns8pGrdeKzh6unEUB64U6gy4RCf4VKa8iJFp7eTldE6pVTJhM5NWZAVdl6L
Arb2jMrv7Pp8szWp6YIXGIRsVchvNw7FRq6IR3U4LM0xCu6rEYI2C4FOawMEmU0f
AUnXZEObBDrkCCl6XZdMqnxszB7ABv0crgGHP/Tq5LnD0Lu38//7PhN0NocpOIm5
liiXsXOpMCanjFeR0mUnAag5W4TGjtNVtSm5IT0KurDE1vNWLK4OpqgKHLGcvviy
wFaSIq2N0rY61RMg0ecFx6zP9iuVa7XZJ8gqmPU4PWOgYIFXI/oUI16XzD6o0Obd
GtaqqoVhT3elYF2sAdek4IcQ6AwBGvBv2Pt6aNzOpTN8SgRgB/2lVBHsjEY2VZv1
PQEvUT3ANhbQMUfqOELuO09J3R4if4Xh8mKz79lcs5+HDaPWxFxI280oXJD6F0iC
JnF8Oph8Q3slBpuB2rHFLfEqPesyr0Br0Z41ljehHIsEgZwJ/A/zXkfzsecwr5NO
GXL3dSkrA6CuGlfFVdbIvDrEfnZZ5ApPci2XJN6iJfbdXb3xHCgfy+ojhX3rit0z
YklFieG+j71sw7mKfclY29bhgS6ts1PyNxWEM42nEqQAuBCcXoz8U1k4f8gvQbRi
klxlWuPA1gnrZ0D1fY1wxLfFQyOrtNo2OhalZmsZuCweFhnH6MJxaJvyyjdtnciS
bvE2fQRuk62tQ3ztO/gWRywvmnn1egw3kuz1ybOEc/Ar+mEoSQNQ1CS5/P5yXTET
k3Zj88lPnwek+XUdTq6FUEnLdM6FrWYLO589VSkrFefSZChcehsbT6vJfF5bQrwq
Fk2VSyyJ/3S11TSG5v5TyC6xv8yifUm3K9ls+LOLrHIMBBkKesXa1lt0Lg580uwF
CaEbfapwkmOZVb7uiK2QbdSGWlKuV7txMIrgh1exgip9Kg4ltDHme4FA80SJnudT
7FsPV92o/UXqUhDREefI8TxMMCyGgs/VrtnV/72WXjYJTWDK3hrHVTruPJWFEhWq
XzHHThVmJ3UiLTIPUMACCg==
`protect END_PROTECTED
